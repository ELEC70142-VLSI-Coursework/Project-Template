VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO PLL_25M_400M
  CLASS BLOCK ;
  ORIGIN -28.225 403.65 ;
  FOREIGN PLL_25M_400M 28.225 -403.65 ;
  SIZE 286.8 BY 194 ;
  SYMMETRY X Y R90 ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M3 ;
        RECT 152.665 -209.975 154.665 -209.65 ;
    END
  END DVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M3 ;
        RECT 157.665 -210.035 159.665 -209.65 ;
    END
    PORT
      LAYER M4 ;
        RECT 267.805 -210.145 269.805 -209.65 ;
    END
  END VSS
  PIN div_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.665 -209.75 182.765 -209.65 ;
    END
  END div_sel[0]
  PIN div_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.665 -209.75 177.765 -209.65 ;
    END
  END div_sel[1]
  PIN div_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.665 -209.75 172.765 -209.65 ;
    END
  END div_sel[2]
  PIN div_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.665 -209.75 167.765 -209.65 ;
    END
  END div_sel[3]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.665 -209.75 162.765 -209.65 ;
    END
  END reset
  PIN CP_20u_Bias
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 272.46 -209.805 272.84 -209.65 ;
    END
  END CP_20u_Bias
  PIN CP_OP_1u_bias
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 273.34 -209.81 273.72 -209.65 ;
    END
  END CP_OP_1u_bias
  PIN f_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.785 -403.65 205.885 -403.55 ;
    END
  END f_out
  PIN input_clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 257.57 -209.75 257.82 -209.65 ;
    END
  END input_clk
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 251.49 -210.18 254.49 -209.65 ;
    END
  END VDD
  OBS
    LAYER M1 SPACING 0.09 ;
      RECT 28.225 -403.65 315.025 -209.65 ;
    LAYER M2 ;
      RECT 273.34 -238.54 273.72 -211.31 ;
      RECT 272.46 -242.71 272.84 -211.305 ;
      RECT 257.57 -212.765 257.82 -211.25 ;
      RECT 205.785 -402.05 206.165 -219.97 ;
    LAYER M2 SPACING 0.1 ;
      RECT 273.91 -403.65 315.025 -209.65 ;
      RECT 273.03 -403.65 273.15 -209.65 ;
      RECT 258.01 -403.65 272.27 -209.65 ;
      RECT 28.225 -403.36 257.38 -209.65 ;
      RECT 28.225 -403.36 272.27 -209.94 ;
      RECT 28.225 -403.36 273.15 -209.995 ;
      RECT 206.075 -403.65 315.025 -210 ;
      RECT 28.225 -403.65 205.595 -209.65 ;
    LAYER M3 ;
      RECT 241.275 -276.8 314.815 -274.83 ;
      RECT 314.395 -319.365 314.815 -274.83 ;
      RECT 184.265 -211.65 184.665 -209.65 ;
      RECT 182.665 -211.65 184.665 -211.25 ;
      RECT 179.265 -211.65 179.665 -209.65 ;
      RECT 177.665 -211.65 179.665 -211.25 ;
      RECT 174.265 -211.65 174.665 -209.65 ;
      RECT 172.665 -211.65 174.665 -211.25 ;
      RECT 169.265 -211.65 169.665 -209.65 ;
      RECT 167.665 -211.65 169.665 -211.25 ;
      RECT 164.265 -211.65 164.665 -209.65 ;
      RECT 162.665 -211.65 164.665 -211.25 ;
      RECT 157.665 -211.65 159.665 -211.535 ;
      RECT 157.715 -215.4 157.815 -211.535 ;
      RECT 152.665 -211.65 154.665 -211.475 ;
      RECT 152.715 -212.4 152.815 -211.475 ;
      RECT 80.955 -378.965 314.815 -372.305 ;
      RECT 80.955 -354.835 314.815 -348.175 ;
    LAYER M3 SPACING 0.1 ;
      RECT 273.91 -403.65 315.025 -209.65 ;
      RECT 273.03 -403.65 273.15 -209.65 ;
      RECT 258.01 -403.65 272.27 -209.65 ;
      RECT 182.955 -403.36 257.38 -209.65 ;
      RECT 177.955 -403.65 182.475 -209.65 ;
      RECT 172.955 -403.65 177.475 -209.65 ;
      RECT 167.955 -403.65 172.475 -209.65 ;
      RECT 162.955 -403.65 167.475 -209.65 ;
      RECT 159.855 -403.65 162.475 -209.65 ;
      RECT 154.855 -403.65 157.475 -209.65 ;
      RECT 28.225 -403.65 152.475 -209.65 ;
      RECT 159.855 -403.36 272.27 -209.94 ;
      RECT 159.855 -403.36 273.15 -209.995 ;
      RECT 206.075 -403.65 315.025 -210 ;
      RECT 28.225 -403.65 157.475 -210.165 ;
      RECT 28.225 -403.65 205.595 -210.225 ;
    LAYER M4 ;
      RECT 28.435 -247.7 87.215 -241.04 ;
      RECT 28.435 -392.01 28.855 -241.04 ;
      RECT 28.435 -272.81 87.215 -266.15 ;
      RECT 28.435 -307.3 262.345 -300.64 ;
      RECT 28.435 -332.41 262.345 -325.75 ;
      RECT 28.435 -366.9 262.345 -360.24 ;
      RECT 28.435 -392.01 262.345 -385.35 ;
      RECT 314.395 -378.965 314.815 -372.305 ;
      RECT 314.395 -354.835 314.815 -348.175 ;
      RECT 314.395 -319.365 314.815 -312.705 ;
      RECT 314.395 -295.235 314.815 -288.575 ;
      RECT 267.805 -243.835 269.805 -211.645 ;
    LAYER M4 SPACING 0.1 ;
      RECT 269.995 -403.65 315.025 -209.65 ;
      RECT 182.955 -403.65 267.615 -209.65 ;
      RECT 177.955 -403.65 182.475 -209.65 ;
      RECT 172.955 -403.65 177.475 -209.65 ;
      RECT 167.955 -403.65 172.475 -209.65 ;
      RECT 162.955 -403.65 167.475 -209.65 ;
      RECT 159.855 -403.65 162.475 -209.65 ;
      RECT 154.855 -403.65 157.475 -209.65 ;
      RECT 28.225 -403.65 152.475 -209.65 ;
      RECT 159.855 -403.65 267.615 -209.94 ;
      RECT 28.225 -403.65 157.475 -210.165 ;
      RECT 28.225 -403.65 267.615 -210.225 ;
      RECT 28.225 -403.65 315.025 -210.335 ;
    LAYER M5 ;
      RECT 314.395 -378.965 314.815 -372.305 ;
      RECT 314.395 -354.835 314.815 -348.175 ;
      RECT 314.395 -319.365 314.815 -312.705 ;
      RECT 314.395 -295.235 314.815 -288.575 ;
      RECT 251.49 -223.355 254.49 -211.68 ;
      RECT 28.435 -392.01 28.855 -385.35 ;
      RECT 28.435 -366.9 28.855 -360.24 ;
      RECT 28.435 -332.41 28.855 -325.75 ;
      RECT 28.435 -307.3 28.855 -300.64 ;
      RECT 28.435 -272.81 28.855 -266.15 ;
      RECT 28.435 -247.7 28.855 -241.04 ;
    LAYER M5 SPACING 0.1 ;
      RECT 269.995 -403.65 315.025 -209.65 ;
      RECT 254.68 -403.65 267.615 -209.65 ;
      RECT 28.225 -403.65 251.3 -209.65 ;
      RECT 254.68 -403.65 315.025 -210.335 ;
      RECT 28.225 -403.65 315.025 -210.37 ;
    LAYER M6 ;
      RECT 314.395 -378.965 314.815 -372.305 ;
      RECT 314.395 -354.835 314.815 -348.175 ;
      RECT 314.395 -319.365 314.815 -312.705 ;
      RECT 314.395 -295.235 314.815 -288.575 ;
      RECT 298.005 -229.95 314.785 -229.55 ;
      RECT 28.435 -392.01 28.855 -385.35 ;
      RECT 28.435 -366.9 28.855 -360.24 ;
      RECT 28.435 -332.41 28.855 -325.75 ;
      RECT 28.435 -307.3 28.855 -300.64 ;
      RECT 28.435 -272.81 28.855 -266.15 ;
      RECT 28.435 -247.7 28.855 -241.04 ;
    LAYER M6 SPACING 0.1 ;
      RECT 254.68 -403.65 315.025 -209.65 ;
      RECT 28.225 -403.65 251.3 -209.65 ;
      RECT 28.225 -403.65 315.025 -210.37 ;
    LAYER M7 ;
      RECT 314.245 -228.25 314.965 -219.85 ;
      RECT 314.405 -251.05 314.805 -219.85 ;
      RECT 314.245 -239.65 314.965 -231.25 ;
      RECT 314.245 -251.05 314.965 -242.65 ;
      RECT 314.345 -379.045 314.865 -372.225 ;
      RECT 314.345 -354.915 314.865 -348.095 ;
      RECT 314.345 -319.445 314.865 -312.625 ;
      RECT 314.345 -295.315 314.865 -288.495 ;
      RECT 28.385 -392.09 28.905 -385.27 ;
      RECT 28.385 -366.98 28.905 -360.16 ;
      RECT 28.385 -332.49 28.905 -325.67 ;
      RECT 28.385 -307.38 28.905 -300.56 ;
      RECT 28.385 -272.89 28.905 -266.07 ;
      RECT 28.385 -247.78 28.905 -240.96 ;
    LAYER M7 SPACING 0.1 ;
      RECT 28.225 -403.65 315.025 -209.65 ;
    LAYER M8 ;
      RECT 263.345 -342.85 315.025 -341.39 ;
      RECT 314.185 -391.11 315.025 -341.39 ;
      RECT 263.345 -354.915 315.025 -353.455 ;
      RECT 263.345 -366.98 315.025 -365.52 ;
      RECT 263.345 -379.045 315.025 -377.585 ;
      RECT 263.345 -391.11 315.025 -389.65 ;
      RECT 263.345 -283.25 315.025 -281.79 ;
      RECT 314.185 -331.51 315.025 -281.79 ;
      RECT 263.345 -295.315 315.025 -293.855 ;
      RECT 263.345 -307.38 315.025 -305.92 ;
      RECT 263.345 -319.445 315.025 -317.985 ;
      RECT 263.345 -331.51 315.025 -330.05 ;
      RECT 313.345 -244.01 315.025 -242.55 ;
      RECT 314.185 -251.15 315.025 -242.55 ;
      RECT 313.345 -251.15 315.025 -249.69 ;
      RECT 313.345 -232.61 315.025 -231.15 ;
      RECT 314.185 -239.75 315.025 -231.15 ;
      RECT 313.345 -239.75 315.025 -238.29 ;
      RECT 313.345 -221.21 315.025 -219.75 ;
      RECT 314.185 -228.35 315.025 -219.75 ;
      RECT 313.345 -228.35 315.025 -226.89 ;
      RECT 28.225 -340.41 29.905 -338.95 ;
      RECT 28.225 -393.55 29.065 -338.95 ;
      RECT 28.225 -393.55 29.905 -392.09 ;
      RECT 28.225 -280.81 29.905 -279.35 ;
      RECT 28.225 -333.95 29.065 -279.35 ;
      RECT 28.225 -333.95 29.905 -332.49 ;
      RECT 28.225 -221.21 29.905 -219.75 ;
      RECT 28.225 -274.35 29.065 -219.75 ;
      RECT 28.225 -274.35 29.905 -272.89 ;
    LAYER M8 SPACING 0.4 ;
      RECT 28.225 -403.65 315.025 -209.65 ;
    LAYER M9 SPACING 2 ;
      RECT 28.225 -403.65 315.025 -209.65 ;
  END
END PLL_25M_400M

END LIBRARY
