* SPICE NETLIST
***************************************

.SUBCKT LDDP D G S B
.ENDS
***************************************
.SUBCKT LDDN D G S B
.ENDS
***************************************
.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_2t PLUS MINUS
.ENDS
***************************************
.SUBCKT crtmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT crtmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT fmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT fmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lincap PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT lincap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lincap_rf_25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT lowcpad_d15 APAD AVSS
.ENDS
***************************************
.SUBCKT lowcpad_d23 APAD AVSS
.ENDS
***************************************
.SUBCKT mimcap_sin PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_um_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_woum_sin_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf18_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf25_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_hvt_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT ndio_hia_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_18_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwod D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25_nodnwud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25od33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_25ud18_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_33_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_cas_nw D GB S B GT
.ENDS
***************************************
.SUBCKT nmos_rf_cross_nw DP DM S B
.ENDS
***************************************
.SUBCKT nmos_rf_diff_nw DP GP S B DM GM
.ENDS
***************************************
.SUBCKT nmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_hvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_lvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_mlvt_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_na18 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_nodnw D G S B
.ENDS
***************************************
.SUBCKT nmos_rf_rdk D G S B
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_18 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_25 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_lpg PLUS MINUS
.ENDS
***************************************
.SUBCKT pdio_hia_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwod D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25_nwud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25od33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_25ud18_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_hvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_lvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_mlvt_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_rdk D G S B
.ENDS
***************************************
.SUBCKT pmoscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf18 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmoscap_rf25 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT probe1 TOP BULK
.ENDS
***************************************
.SUBCKT probe2 TOP BULK
.ENDS
***************************************
.SUBCKT probe3 TOP BULK
.ENDS
***************************************
.SUBCKT probe4 TOP BULK
.ENDS
***************************************
.SUBCKT probe5 TOP BULK
.ENDS
***************************************
.SUBCKT probe6 TOP BULK
.ENDS
***************************************
.SUBCKT probe7 TOP BULK
.ENDS
***************************************
.SUBCKT rfesd_rf1 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf2 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf3 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf4 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf5 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf6 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf7 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rfesd_rf8 APAD CPAD DCPAD GNODE
.ENDS
***************************************
.SUBCKT rm1 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm10 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm2 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm3 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm4 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm5 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm6 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm7 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm8 PLUS MINUS
.ENDS
***************************************
.SUBCKT rm9 PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnods PLUS MINUS
.ENDS
***************************************
.SUBCKT rnods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnpolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwod PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rnwsti PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodl PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpods PLUS MINUS
.ENDS
***************************************
.SUBCKT rpods_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rpodwo PLUS MINUS
.ENDS
***************************************
.SUBCKT rpodwo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolyl_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolys_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo PLUS MINUS
.ENDS
***************************************
.SUBCKT rppolywo_m PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sline_gscpw_mu PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sline_ms_mu PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_z_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_z_rdk PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_mu_z_rdk PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_CDNS_764966941090 1 2
** N=2 EP=2 IP=0 FDC=1
X0 2 1 mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=0 $Y=0 $D=325
.ENDS
***************************************
.SUBCKT FILL2BWP7T
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILL1BWP7T
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_5
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT DCAP16BWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=8
M0 VSS 3 VSS VSS nch L=6.25e-07 W=1.7e-07 $X=225 $Y=260 $D=4
M1 VSS 3 VSS VSS nch L=6.1e-07 W=1.7e-07 $X=1150 $Y=260 $D=4
M2 VSS 3 VSS VSS nch L=6.1e-07 W=1.7e-07 $X=2035 $Y=260 $D=4
M3 4 3 VSS VSS nch L=6e-08 W=1.7e-07 $X=2915 $Y=260 $D=4
M4 VDD 4 VDD VDD pch L=6.1e-07 W=2.15e-07 $X=240 $Y=925 $D=103
M5 VDD 4 VDD VDD pch L=6.1e-07 W=2.15e-07 $X=1150 $Y=925 $D=103
M6 VDD 4 VDD VDD pch L=6.1e-07 W=2.15e-07 $X=2035 $Y=925 $D=103
M7 3 4 VDD VDD pch L=6e-08 W=2.15e-07 $X=2850 $Y=925 $D=103
.ENDS
***************************************
.SUBCKT ICV_11 1 2
** N=2 EP=2 IP=4 FDC=8
X1 2 1 DCAP16BWP7T $T=0 0 0 0 $X=-235 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_17 1 2
** N=2 EP=2 IP=4 FDC=8
X1 1 2 ICV_11 $T=600 0 0 0 $X=365 $Y=-105
.ENDS
***************************************
.SUBCKT DCAP4BWP7T VSS VDD
** N=4 EP=2 IP=0 FDC=4
M0 VSS 4 VSS VSS nch L=6e-08 W=2.5e-07 $X=240 $Y=200 $D=4
M1 3 4 VSS VSS nch L=6e-08 W=2.5e-07 $X=505 $Y=200 $D=4
M2 VDD 3 VDD VDD pch L=6e-08 W=3.2e-07 $X=250 $Y=880 $D=103
M3 4 3 VDD VDD pch L=6e-08 W=3.2e-07 $X=515 $Y=880 $D=103
.ENDS
***************************************
.SUBCKT TAPCELLBWP7T
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_9 1 2
** N=2 EP=2 IP=4 FDC=4
X0 1 2 DCAP4BWP7T $T=0 0 0 0 $X=-235 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_18 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 ICV_9 $T=0 0 0 0 $X=-235 $Y=-105
.ENDS
***************************************
.SUBCKT DCAP32BWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=16
M0 VSS 3 4 VSS nch L=6e-08 W=1.7e-07 $X=230 $Y=260 $D=4
M1 VSS 3 VSS VSS nch L=6e-07 W=1.7e-07 $X=570 $Y=260 $D=4
M2 VSS 3 VSS VSS nch L=6.1e-07 W=1.7e-07 $X=1445 $Y=260 $D=4
M3 VSS 3 VSS VSS nch L=6.95e-07 W=1.7e-07 $X=2355 $Y=260 $D=4
M4 VSS 3 VSS VSS nch L=6.6e-07 W=1.7e-07 $X=3390 $Y=260 $D=4
M5 VSS 3 VSS VSS nch L=6.1e-07 W=1.7e-07 $X=4350 $Y=260 $D=4
M6 VSS 3 VSS VSS nch L=5.95e-07 W=1.7e-07 $X=5235 $Y=260 $D=4
M7 4 3 VSS VSS nch L=6e-08 W=1.7e-07 $X=6115 $Y=260 $D=4
M8 VDD 4 3 VDD pch L=6e-08 W=2.15e-07 $X=295 $Y=925 $D=103
M9 VDD 4 VDD VDD pch L=6.1e-07 W=2.15e-07 $X=560 $Y=925 $D=103
M10 VDD 4 VDD VDD pch L=6.1e-07 W=2.15e-07 $X=1445 $Y=925 $D=103
M11 VDD 4 VDD VDD pch L=6.95e-07 W=2.15e-07 $X=2355 $Y=925 $D=103
M12 VDD 4 VDD VDD pch L=6.6e-07 W=2.15e-07 $X=3390 $Y=925 $D=103
M13 VDD 4 VDD VDD pch L=6.1e-07 W=2.15e-07 $X=4350 $Y=925 $D=103
M14 VDD 4 VDD VDD pch L=6.1e-07 W=2.15e-07 $X=5235 $Y=925 $D=103
M15 3 4 VDD VDD pch L=6e-08 W=2.15e-07 $X=6050 $Y=925 $D=103
.ENDS
***************************************
.SUBCKT DCAP8BWP7T VDD VSS
** N=4 EP=2 IP=0 FDC=4
M0 VSS 3 VSS VSS nch L=8.05e-07 W=1.7e-07 $X=225 $Y=260 $D=4
M1 4 3 VSS VSS nch L=6e-08 W=1.7e-07 $X=1315 $Y=260 $D=4
M2 VDD 4 VDD VDD pch L=8.1e-07 W=2.2e-07 $X=240 $Y=920 $D=103
M3 3 4 VDD VDD pch L=6e-08 W=2.2e-07 $X=1250 $Y=920 $D=103
.ENDS
***************************************
.SUBCKT ICV_1 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 DCAP4BWP7T $T=200 0 0 0 $X=-35 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_12 1 2
** N=2 EP=2 IP=6 FDC=24
X0 1 2 DCAP32BWP7T $T=0 0 0 0 $X=-235 $Y=-105
X1 1 2 DCAP8BWP7T $T=6400 0 0 0 $X=6165 $Y=-105
X2 2 1 ICV_1 $T=8000 0 0 0 $X=7765 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_19 1 2
** N=2 EP=2 IP=12 FDC=72
X0 1 2 ICV_17 $T=0 0 0 0 $X=-235 $Y=-105
X1 1 2 ICV_17 $T=0 2800 1 0 $X=-235 $Y=1165
X2 1 2 ICV_18 $T=4200 0 0 0 $X=3965 $Y=-105
X3 1 2 ICV_18 $T=4200 2800 1 0 $X=3965 $Y=1165
X4 2 1 ICV_12 $T=6000 0 0 0 $X=5765 $Y=-105
X5 2 1 ICV_12 $T=6000 2800 1 0 $X=5765 $Y=1165
.ENDS
***************************************
.SUBCKT ICV_4 1 2
** N=2 EP=2 IP=4 FDC=4
X1 2 1 DCAP8BWP7T $T=0 0 0 0 $X=-235 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_13 1 2
** N=2 EP=2 IP=4 FDC=4
X1 1 2 ICV_1 $T=600 0 0 0 $X=365 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_10 1 2
** N=2 EP=2 IP=4 FDC=4
X1 2 1 DCAP8BWP7T $T=200 0 0 0 $X=-35 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_14
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15 1 2
** N=2 EP=2 IP=6 FDC=20
X0 1 2 DCAP32BWP7T $T=0 0 0 0 $X=-235 $Y=-105
X1 2 1 ICV_10 $T=6400 0 0 0 $X=6165 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_16 1 2
** N=2 EP=2 IP=14 FDC=44
X3 2 1 DCAP32BWP7T $T=1800 0 0 0 $X=1565 $Y=-105
X4 1 2 ICV_4 $T=8200 0 0 0 $X=7965 $Y=-105
X5 1 2 ICV_13 $T=0 0 0 0 $X=-235 $Y=-105
X6 2 1 ICV_15 $T=11200 0 0 0 $X=10965 $Y=-105
.ENDS
***************************************
.SUBCKT FILL32BWP7T
** N=51 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILL8BWP7T
** N=12 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILL16BWP7T
** N=27 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2 1 2
** N=2 EP=2 IP=4 FDC=8
X1 2 1 DCAP16BWP7T $T=200 0 0 0 $X=-35 $Y=-105
.ENDS
***************************************
.SUBCKT DFKCNQD1BWP7T CP CN D VDD VSS Q
** N=18 EP=6 IP=0 FDC=26
M0 VSS CP 9 VSS nch L=6e-08 W=1.5e-07 $X=225 $Y=350 $D=4
M1 11 9 VSS VSS nch L=6e-08 W=1.5e-07 $X=470 $Y=350 $D=4
M2 16 CN VSS VSS nch L=6e-08 W=2.8e-07 $X=950 $Y=220 $D=4
M3 17 D 16 VSS nch L=6e-08 W=2.8e-07 $X=1185 $Y=220 $D=4
M4 8 9 17 VSS nch L=6e-08 W=2.8e-07 $X=1420 $Y=220 $D=4
M5 18 11 8 VSS nch L=6e-08 W=1.5e-07 $X=1845 $Y=350 $D=4
M6 VSS 10 18 VSS nch L=6e-08 W=1.5e-07 $X=2095 $Y=350 $D=4
M7 10 8 VSS VSS nch L=6e-08 W=2.7e-07 $X=2405 $Y=265 $D=4
M8 12 11 10 VSS nch L=6e-08 W=1.5e-07 $X=2690 $Y=350 $D=4
M9 13 9 12 VSS nch L=6e-08 W=1.5e-07 $X=3045 $Y=250 $D=4
M10 VSS 14 13 VSS nch L=6e-08 W=1.5e-07 $X=3385 $Y=250 $D=4
M11 14 12 VSS VSS nch L=6e-08 W=1.9e-07 $X=3635 $Y=345 $D=4
M12 Q 14 VSS VSS nch L=6e-08 W=2.8e-07 $X=4110 $Y=220 $D=4
M13 VDD CP 9 VDD pch L=6e-08 W=1.9e-07 $X=225 $Y=820 $D=103
M14 11 9 VDD VDD pch L=6e-08 W=1.9e-07 $X=470 $Y=820 $D=103
M15 VDD CN 7 VDD pch L=6e-08 W=1.9e-07 $X=960 $Y=820 $D=103
M16 7 D VDD VDD pch L=6e-08 W=3.6e-07 $X=1200 $Y=820 $D=103
M17 8 11 7 VDD pch L=6e-08 W=1.95e-07 $X=1545 $Y=985 $D=103
M18 15 9 8 VDD pch L=6e-08 W=1.5e-07 $X=1930 $Y=900 $D=103
M19 VDD 10 15 VDD pch L=6e-08 W=1.5e-07 $X=2155 $Y=900 $D=103
M20 10 8 VDD VDD pch L=6e-08 W=3.25e-07 $X=2475 $Y=855 $D=103
M21 12 9 10 VDD pch L=6e-08 W=1.5e-07 $X=2820 $Y=900 $D=103
M22 13 11 12 VDD pch L=6e-08 W=1.5e-07 $X=3095 $Y=900 $D=103
M23 VDD 14 13 VDD pch L=6e-08 W=1.9e-07 $X=3385 $Y=900 $D=103
M24 14 12 VDD VDD pch L=6e-08 W=1.9e-07 $X=3635 $Y=855 $D=103
M25 Q 14 VDD VDD pch L=6e-08 W=3.25e-07 $X=4110 $Y=855 $D=103
.ENDS
***************************************
.SUBCKT FILL4BWP7T
** N=6 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT HA1D0BWP7T CO B A VSS VDD S
** N=13 EP=6 IP=0 FDC=18
M0 VSS 7 CO VSS nch L=6e-08 W=1.5e-07 $X=215 $Y=200 $D=4
M1 12 B VSS VSS nch L=6e-08 W=1.5e-07 $X=485 $Y=380 $D=4
M2 7 A 12 VSS nch L=6e-08 W=1.5e-07 $X=685 $Y=380 $D=4
M3 VSS A 8 VSS nch L=6e-08 W=1.5e-07 $X=1175 $Y=380 $D=4
M4 13 8 VSS VSS nch L=6e-08 W=1.5e-07 $X=1435 $Y=380 $D=4
M5 10 B 13 VSS nch L=6e-08 W=1.5e-07 $X=1625 $Y=380 $D=4
M6 8 9 10 VSS nch L=6e-08 W=1.5e-07 $X=1895 $Y=380 $D=4
M7 VSS B 9 VSS nch L=6e-08 W=1.5e-07 $X=2465 $Y=275 $D=4
M8 S 10 VSS VSS nch L=6e-08 W=1.5e-07 $X=2725 $Y=275 $D=4
M9 VDD 7 CO VDD pch L=6e-08 W=1.9e-07 $X=215 $Y=850 $D=103
M10 7 B VDD VDD pch L=6e-08 W=1.9e-07 $X=455 $Y=850 $D=103
M11 VDD A 7 VDD pch L=6e-08 W=1.9e-07 $X=715 $Y=850 $D=103
M12 VDD A 8 VDD pch L=6e-08 W=2.65e-07 $X=1195 $Y=915 $D=103
M13 11 8 VDD VDD pch L=6e-08 W=2.3e-07 $X=1455 $Y=970 $D=103
M14 10 9 11 VDD pch L=6e-08 W=2.3e-07 $X=1670 $Y=970 $D=103
M15 8 B 10 VDD pch L=6e-08 W=1.9e-07 $X=1985 $Y=1010 $D=103
M16 VDD B 9 VDD pch L=6e-08 W=1.9e-07 $X=2485 $Y=820 $D=103
M17 S 10 VDD VDD pch L=6e-08 W=1.9e-07 $X=2725 $Y=820 $D=103
.ENDS
***************************************
.SUBCKT OAI31D1BWP7T A1 A2 A3 ZN B VDD VSS
** N=10 EP=7 IP=0 FDC=8
M0 8 A1 ZN VSS nch L=6e-08 W=3e-07 $X=225 $Y=200 $D=4
M1 ZN A2 8 VSS nch L=6e-08 W=3e-07 $X=490 $Y=200 $D=4
M2 8 A3 ZN VSS nch L=6e-08 W=3e-07 $X=755 $Y=200 $D=4
M3 VSS B 8 VSS nch L=6e-08 W=3e-07 $X=1065 $Y=200 $D=4
M4 9 A1 VDD VDD pch L=6e-08 W=3.8e-07 $X=225 $Y=820 $D=103
M5 10 A2 9 VDD pch L=6e-08 W=3.8e-07 $X=490 $Y=820 $D=103
M6 ZN A3 10 VDD pch L=6e-08 W=3.8e-07 $X=755 $Y=820 $D=103
M7 VDD B ZN VDD pch L=6e-08 W=3.8e-07 $X=1065 $Y=820 $D=103
.ENDS
***************************************
.SUBCKT AOI21D0BWP7T A2 ZN A1 B VDD VSS
** N=8 EP=6 IP=0 FDC=6
M0 8 A2 VSS VSS nch L=6e-08 W=1.5e-07 $X=215 $Y=200 $D=4
M1 ZN A1 8 VSS nch L=6e-08 W=1.5e-07 $X=415 $Y=200 $D=4
M2 VSS B ZN VSS nch L=6e-08 W=1.5e-07 $X=695 $Y=200 $D=4
M3 ZN A2 7 VDD pch L=6e-08 W=1.9e-07 $X=195 $Y=860 $D=103
M4 7 A1 ZN VDD pch L=6e-08 W=1.9e-07 $X=455 $Y=860 $D=103
M5 VDD B 7 VDD pch L=6e-08 W=1.9e-07 $X=695 $Y=860 $D=103
.ENDS
***************************************
.SUBCKT MUX2ND0BWP7T I0 S ZN I1 VSS VDD
** N=11 EP=6 IP=0 FDC=10
M0 VSS S 7 VSS nch L=6e-08 W=1.5e-07 $X=225 $Y=200 $D=4
M1 10 I0 VSS VSS nch L=6e-08 W=1.5e-07 $X=485 $Y=200 $D=4
M2 ZN 7 10 VSS nch L=6e-08 W=1.5e-07 $X=710 $Y=200 $D=4
M3 11 S ZN VSS nch L=6e-08 W=1.5e-07 $X=975 $Y=200 $D=4
M4 VSS I1 11 VSS nch L=6e-08 W=1.5e-07 $X=1265 $Y=200 $D=4
M5 VDD S 7 VDD pch L=6e-08 W=1.9e-07 $X=225 $Y=820 $D=103
M6 8 I0 VDD VDD pch L=6e-08 W=1.8e-07 $X=505 $Y=820 $D=103
M7 ZN S 8 VDD pch L=6e-08 W=1.9e-07 $X=765 $Y=1010 $D=103
M8 9 7 ZN VDD pch L=6e-08 W=1.9e-07 $X=1040 $Y=1010 $D=103
M9 VDD I1 9 VDD pch L=6e-08 W=1.9e-07 $X=1265 $Y=1010 $D=103
.ENDS
***************************************
.SUBCKT ICV_8
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT IND2D1BWP7T A1 VSS ZN B1 VDD
** N=7 EP=5 IP=0 FDC=6
M0 VSS A1 6 VSS nch L=6e-08 W=1.5e-07 $X=215 $Y=200 $D=4
M1 7 6 VSS VSS nch L=6e-08 W=3e-07 $X=475 $Y=200 $D=4
M2 ZN B1 7 VSS nch L=6e-08 W=3e-07 $X=705 $Y=200 $D=4
M3 VDD A1 6 VDD pch L=6e-08 W=1.9e-07 $X=215 $Y=820 $D=103
M4 ZN 6 VDD VDD pch L=6e-08 W=3.6e-07 $X=455 $Y=820 $D=103
M5 VDD B1 ZN VDD pch L=6e-08 W=3.8e-07 $X=715 $Y=820 $D=103
.ENDS
***************************************
.SUBCKT IOA21D0BWP7T A1 A2 VSS ZN B VDD
** N=9 EP=6 IP=0 FDC=8
M0 8 A1 7 VSS nch L=6e-08 W=1.5e-07 $X=215 $Y=220 $D=4
M1 VSS A2 8 VSS nch L=6e-08 W=1.5e-07 $X=415 $Y=220 $D=4
M2 9 7 VSS VSS nch L=6e-08 W=1.5e-07 $X=725 $Y=220 $D=4
M3 ZN B 9 VSS nch L=6e-08 W=1.5e-07 $X=925 $Y=220 $D=4
M4 7 A1 VDD VDD pch L=6e-08 W=1.8e-07 $X=190 $Y=835 $D=103
M5 VDD A2 7 VDD pch L=6e-08 W=1.8e-07 $X=450 $Y=835 $D=103
M6 ZN 7 VDD VDD pch L=6e-08 W=1.8e-07 $X=690 $Y=835 $D=103
M7 VDD B ZN VDD pch L=6e-08 W=1.8e-07 $X=950 $Y=835 $D=103
.ENDS
***************************************
.SUBCKT EDFKCNQD1BWP7T E D CN CP VSS VDD Q
** N=23 EP=7 IP=0 FDC=34
M0 8 E VSS VSS nch L=6e-08 W=1.5e-07 $X=235 $Y=350 $D=4
M1 21 17 9 VSS nch L=6e-08 W=1.5e-07 $X=725 $Y=380 $D=4
M2 12 8 21 VSS nch L=6e-08 W=1.5e-07 $X=925 $Y=380 $D=4
M3 22 E 12 VSS nch L=6e-08 W=2.3e-07 $X=1200 $Y=200 $D=4
M4 9 D 22 VSS nch L=6e-08 W=2.3e-07 $X=1400 $Y=200 $D=4
M5 VSS CN 9 VSS nch L=6e-08 W=2.3e-07 $X=1660 $Y=200 $D=4
M6 VSS CP 10 VSS nch L=6e-08 W=1.5e-07 $X=2255 $Y=385 $D=4
M7 11 10 VSS VSS nch L=6e-08 W=1.5e-07 $X=2495 $Y=385 $D=4
M8 13 10 12 VSS nch L=6e-08 W=1.5e-07 $X=3010 $Y=200 $D=4
M9 23 11 13 VSS nch L=6e-08 W=1.5e-07 $X=3290 $Y=220 $D=4
M10 VSS 14 23 VSS nch L=6e-08 W=1.5e-07 $X=3490 $Y=220 $D=4
M11 14 13 VSS VSS nch L=6e-08 W=3.05e-07 $X=3800 $Y=230 $D=4
M12 15 11 14 VSS nch L=6e-08 W=1.5e-07 $X=4135 $Y=350 $D=4
M13 17 10 15 VSS nch L=6e-08 W=1.5e-07 $X=4460 $Y=220 $D=4
M14 VSS 16 17 VSS nch L=6e-08 W=1.5e-07 $X=4800 $Y=220 $D=4
M15 16 15 VSS VSS nch L=6e-08 W=1.9e-07 $X=5040 $Y=345 $D=4
M16 Q 16 VSS VSS nch L=6e-08 W=2.8e-07 $X=5515 $Y=220 $D=4
M17 VDD E 8 VDD pch L=6e-08 W=1.5e-07 $X=225 $Y=895 $D=103
M18 18 E VDD VDD pch L=6e-08 W=1.7e-07 $X=535 $Y=1010 $D=103
M19 12 17 18 VDD pch L=6e-08 W=1.7e-07 $X=760 $Y=1010 $D=103
M20 19 8 12 VDD pch L=6e-08 W=3.5e-07 $X=1100 $Y=850 $D=103
M21 VDD D 19 VDD pch L=6e-08 W=3.5e-07 $X=1300 $Y=850 $D=103
M22 12 CN VDD VDD pch L=6e-08 W=1.5e-07 $X=1710 $Y=850 $D=103
M23 VDD CP 10 VDD pch L=6e-08 W=1.9e-07 $X=2290 $Y=855 $D=103
M24 11 10 VDD VDD pch L=6e-08 W=1.9e-07 $X=2530 $Y=855 $D=103
M25 13 11 12 VDD pch L=6e-08 W=1.65e-07 $X=3020 $Y=855 $D=103
M26 20 10 13 VDD pch L=6e-08 W=1.5e-07 $X=3300 $Y=950 $D=103
M27 VDD 14 20 VDD pch L=6e-08 W=1.65e-07 $X=3575 $Y=855 $D=103
M28 14 13 VDD VDD pch L=6e-08 W=1.65e-07 $X=3955 $Y=855 $D=103
M29 15 10 14 VDD pch L=6e-08 W=1.5e-07 $X=4265 $Y=900 $D=103
M30 17 11 15 VDD pch L=6e-08 W=1.5e-07 $X=4525 $Y=900 $D=103
M31 VDD 16 17 VDD pch L=6e-08 W=1.5e-07 $X=4825 $Y=900 $D=103
M32 16 15 VDD VDD pch L=6e-08 W=1.9e-07 $X=5065 $Y=865 $D=103
M33 Q 16 VDD VDD pch L=6e-08 W=3.25e-07 $X=5525 $Y=855 $D=103
.ENDS
***************************************
.SUBCKT XOR2D1BWP7T A1 A2 VDD VSS Z
** N=10 EP=5 IP=0 FDC=12
M0 VSS A1 6 VSS nch L=6e-08 W=1.5e-07 $X=215 $Y=350 $D=4
M1 10 7 VSS VSS nch L=6e-08 W=1.5e-07 $X=545 $Y=380 $D=4
M2 8 A1 10 VSS nch L=6e-08 W=1.5e-07 $X=835 $Y=200 $D=4
M3 7 6 8 VSS nch L=6e-08 W=1.5e-07 $X=1095 $Y=200 $D=4
M4 VSS A2 7 VSS nch L=6e-08 W=1.5e-07 $X=1385 $Y=385 $D=4
M5 Z 8 VSS VSS nch L=6e-08 W=2.8e-07 $X=1715 $Y=220 $D=4
M6 VDD A1 6 VDD pch L=6e-08 W=1.9e-07 $X=215 $Y=1010 $D=103
M7 9 7 VDD VDD pch L=6e-08 W=1.5e-07 $X=515 $Y=850 $D=103
M8 8 6 9 VDD pch L=6e-08 W=1.5e-07 $X=725 $Y=850 $D=103
M9 7 A1 8 VDD pch L=6e-08 W=1.9e-07 $X=995 $Y=1010 $D=103
M10 VDD A2 7 VDD pch L=6e-08 W=1.9e-07 $X=1305 $Y=1010 $D=103
M11 Z 8 VDD VDD pch L=6e-08 W=3.45e-07 $X=1715 $Y=855 $D=103
.ENDS
***************************************
.SUBCKT INR2XD0BWP7T A1 VDD ZN B1 VSS
** N=7 EP=5 IP=0 FDC=6
M0 VSS A1 6 VSS nch L=6e-08 W=1.5e-07 $X=215 $Y=350 $D=4
M1 ZN 6 VSS VSS nch L=6e-08 W=1.5e-07 $X=455 $Y=350 $D=4
M2 VSS B1 ZN VSS nch L=6e-08 W=1.5e-07 $X=715 $Y=350 $D=4
M3 VDD A1 6 VDD pch L=6e-08 W=1.9e-07 $X=215 $Y=1010 $D=103
M4 7 6 VDD VDD pch L=6e-08 W=3.8e-07 $X=475 $Y=820 $D=103
M5 ZN B1 7 VDD pch L=6e-08 W=3.8e-07 $X=685 $Y=820 $D=103
.ENDS
***************************************
.SUBCKT XNR2D1BWP7T A1 A2 VDD VSS ZN
** N=10 EP=5 IP=0 FDC=12
M0 VSS A1 6 VSS nch L=6e-08 W=1.5e-07 $X=215 $Y=200 $D=4
M1 10 7 VSS VSS nch L=6e-08 W=1.5e-07 $X=535 $Y=380 $D=4
M2 8 6 10 VSS nch L=6e-08 W=1.5e-07 $X=735 $Y=380 $D=4
M3 7 A1 8 VSS nch L=6e-08 W=1.5e-07 $X=1055 $Y=200 $D=4
M4 VSS A2 7 VSS nch L=6e-08 W=3e-07 $X=1355 $Y=230 $D=4
M5 ZN 8 VSS VSS nch L=6e-08 W=2.8e-07 $X=1715 $Y=220 $D=4
M6 VDD A1 6 VDD pch L=6e-08 W=1.9e-07 $X=215 $Y=1010 $D=103
M7 9 7 VDD VDD pch L=6e-08 W=1.5e-07 $X=500 $Y=850 $D=103
M8 8 A1 9 VDD pch L=6e-08 W=1.7e-07 $X=760 $Y=1030 $D=103
M9 7 6 8 VDD pch L=6e-08 W=1.9e-07 $X=1050 $Y=850 $D=103
M10 VDD A2 7 VDD pch L=6e-08 W=3.5e-07 $X=1355 $Y=850 $D=103
M11 ZN 8 VDD VDD pch L=6e-08 W=3.5e-07 $X=1715 $Y=850 $D=103
.ENDS
***************************************
.SUBCKT BUFFD1BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS I 5 VSS nch L=6e-08 W=1.5e-07 $X=225 $Y=200 $D=4
M1 Z 5 VSS VSS nch L=6e-08 W=3e-07 $X=505 $Y=200 $D=4
M2 VDD I 5 VDD pch L=6e-08 W=1.9e-07 $X=225 $Y=1010 $D=103
M3 Z 5 VDD VDD pch L=6e-08 W=3.8e-07 $X=505 $Y=820 $D=103
.ENDS
***************************************
.SUBCKT ICV_3 1 2
** N=2 EP=2 IP=4 FDC=8
X1 1 2 ICV_2 $T=0 0 0 0 $X=-235 $Y=-105
.ENDS
***************************************
.SUBCKT ICV_7 1 2
** N=2 EP=2 IP=6 FDC=12
X0 1 2 DCAP4BWP7T $T=800 0 0 0 $X=565 $Y=-105
X2 1 2 ICV_3 $T=1600 0 0 0 $X=1365 $Y=-105
.ENDS
***************************************
.SUBCKT clk_div VDD VSS clk_out clk rst_n div_sel[1] div_sel[2] div_sel[3] div_sel[0]
** N=147 EP=9 IP=624 FDC=2248
M0 VSS 10 11 VSS nch L=6e-08 W=3e-07 $X=10250 $Y=10900 $D=4
M1 clk_out 11 VSS VSS nch L=6e-08 W=3e-07 $X=10655 $Y=10900 $D=4
M2 VSS 11 clk_out VSS nch L=6e-08 W=3e-07 $X=10915 $Y=10900 $D=4
M3 VSS 40 12 VSS nch L=6e-08 W=2.8e-07 $X=27030 $Y=13700 $D=4
M4 13 15 VSS VSS nch L=6e-08 W=2.8e-07 $X=27340 $Y=13700 $D=4
M5 VSS 17 15 VSS nch L=6e-08 W=1.9e-07 $X=27890 $Y=13665 $D=4
M6 40 15 VSS VSS nch L=6e-08 W=1.5e-07 $X=28140 $Y=13830 $D=4
M7 17 30 40 VSS nch L=6e-08 W=1.5e-07 $X=28480 $Y=13830 $D=4
M8 18 21 17 VSS nch L=6e-08 W=1.5e-07 $X=28795 $Y=13700 $D=4
M9 VSS 20 10 VSS nch L=6e-08 W=1.5e-07 $X=29015 $Y=11050 $D=4
M10 VSS 22 18 VSS nch L=6e-08 W=3.05e-07 $X=29130 $Y=13665 $D=4
M11 127 19 VSS VSS nch L=6e-08 W=1.5e-07 $X=29275 $Y=11050 $D=4
M12 128 18 VSS VSS nch L=6e-08 W=1.5e-07 $X=29440 $Y=13830 $D=4
M13 20 26 127 VSS nch L=6e-08 W=1.5e-07 $X=29565 $Y=11050 $D=4
M14 22 21 128 VSS nch L=6e-08 W=1.5e-07 $X=29640 $Y=13830 $D=4
M15 129 27 20 VSS nch L=6e-08 W=1.5e-07 $X=29830 $Y=11050 $D=4
M16 39 30 22 VSS nch L=6e-08 W=1.5e-07 $X=29920 $Y=13850 $D=4
M17 VSS clk 129 VSS nch L=6e-08 W=1.5e-07 $X=30055 $Y=11050 $D=4
M18 VSS 37 25 VSS nch L=6e-08 W=2.8e-07 $X=30230 $Y=24900 $D=4
M19 27 26 VSS VSS nch L=6e-08 W=1.5e-07 $X=30315 $Y=11050 $D=4
M20 VSS 30 21 VSS nch L=6e-08 W=1.5e-07 $X=30445 $Y=13665 $D=4
M21 31 36 VSS VSS nch L=6e-08 W=2.8e-07 $X=30540 $Y=24900 $D=4
M22 30 32 VSS VSS nch L=6e-08 W=1.5e-07 $X=30685 $Y=13665 $D=4
M23 VSS 38 36 VSS nch L=6e-08 W=1.9e-07 $X=31105 $Y=24865 $D=4
M24 41 28 VSS VSS nch L=6e-08 W=2.3e-07 $X=31280 $Y=13770 $D=4
M25 37 36 VSS VSS nch L=6e-08 W=1.5e-07 $X=31355 $Y=25000 $D=4
M26 130 12 41 VSS nch L=6e-08 W=2.3e-07 $X=31540 $Y=13770 $D=4
M27 38 48 37 VSS nch L=6e-08 W=1.5e-07 $X=31695 $Y=25000 $D=4
M28 39 47 130 VSS nch L=6e-08 W=2.3e-07 $X=31740 $Y=13770 $D=4
M29 42 46 38 VSS nch L=6e-08 W=1.5e-07 $X=32000 $Y=24900 $D=4
M30 131 43 39 VSS nch L=6e-08 W=1.5e-07 $X=32015 $Y=13670 $D=4
M31 41 40 131 VSS nch L=6e-08 W=1.5e-07 $X=32215 $Y=13670 $D=4
M32 VSS 44 42 VSS nch L=6e-08 W=2.7e-07 $X=32335 $Y=24865 $D=4
M33 132 42 VSS VSS nch L=6e-08 W=1.5e-07 $X=32645 $Y=24900 $D=4
M34 VSS 47 43 VSS nch L=6e-08 W=1.5e-07 $X=32705 $Y=13700 $D=4
M35 44 46 132 VSS nch L=6e-08 W=1.5e-07 $X=32895 $Y=24900 $D=4
M36 133 48 44 VSS nch L=6e-08 W=2.8e-07 $X=33320 $Y=24900 $D=4
M37 134 28 133 VSS nch L=6e-08 W=2.8e-07 $X=33555 $Y=24900 $D=4
M38 VSS 25 134 VSS nch L=6e-08 W=2.8e-07 $X=33790 $Y=24900 $D=4
M39 VSS 48 46 VSS nch L=6e-08 W=1.5e-07 $X=34270 $Y=24900 $D=4
M40 48 32 VSS VSS nch L=6e-08 W=1.5e-07 $X=34515 $Y=24900 $D=4
M41 VSS 50 52 VSS nch L=6e-08 W=1.5e-07 $X=38450 $Y=17200 $D=4
M42 135 49 VSS VSS nch L=6e-08 W=1.5e-07 $X=38710 $Y=17200 $D=4
M43 55 52 135 VSS nch L=6e-08 W=1.5e-07 $X=38910 $Y=17200 $D=4
M44 136 50 55 VSS nch L=6e-08 W=1.5e-07 $X=39175 $Y=17200 $D=4
M45 137 34 VSS VSS nch L=6e-08 W=1.5e-07 $X=39215 $Y=22220 $D=4
M46 138 51 137 VSS nch L=6e-08 W=1.5e-07 $X=39415 $Y=22220 $D=4
M47 VSS 53 136 VSS nch L=6e-08 W=1.5e-07 $X=39435 $Y=17200 $D=4
M48 56 54 138 VSS nch L=6e-08 W=1.5e-07 $X=39690 $Y=22100 $D=4
M49 60 55 VSS VSS nch L=6e-08 W=3e-07 $X=39715 $Y=17200 $D=4
M50 138 60 56 VSS nch L=6e-08 W=1.5e-07 $X=39950 $Y=22100 $D=4
M51 VSS 74 68 VSS nch L=6e-08 W=2.8e-07 $X=46225 $Y=13700 $D=4
M52 69 72 VSS VSS nch L=6e-08 W=2.55e-07 $X=46540 $Y=13700 $D=4
M53 76 68 VSS VSS nch L=6e-08 W=1.5e-07 $X=46820 $Y=17200 $D=4
M54 VSS 75 63 VSS nch L=6e-08 W=2.05e-07 $X=47025 $Y=14400 $D=4
M55 VSS 66 76 VSS nch L=6e-08 W=1.5e-07 $X=47080 $Y=17200 $D=4
M56 VSS 79 72 VSS nch L=6e-08 W=1.9e-07 $X=47105 $Y=13665 $D=4
M57 VSS 26 71 VSS nch L=6e-08 W=1.5e-07 $X=47285 $Y=22800 $D=4
M58 139 69 VSS VSS nch L=6e-08 W=2.05e-07 $X=47295 $Y=14400 $D=4
M59 76 53 VSS VSS nch L=6e-08 W=1.5e-07 $X=47340 $Y=17200 $D=4
M60 74 72 VSS VSS nch L=6e-08 W=1.5e-07 $X=47355 $Y=13830 $D=4
M61 75 77 139 VSS nch L=6e-08 W=2.05e-07 $X=47515 $Y=14400 $D=4
M62 78 71 VSS VSS nch L=6e-08 W=1.5e-07 $X=47595 $Y=22800 $D=4
M63 VSS 65 76 VSS nch L=6e-08 W=1.5e-07 $X=47600 $Y=17200 $D=4
M64 79 91 74 VSS nch L=6e-08 W=1.5e-07 $X=47695 $Y=13830 $D=4
M65 VSS 77 78 VSS nch L=6e-08 W=1.5e-07 $X=47855 $Y=22800 $D=4
M66 26 76 VSS VSS nch L=6e-08 W=3e-07 $X=47860 $Y=17200 $D=4
M67 83 89 79 VSS nch L=6e-08 W=1.5e-07 $X=48000 $Y=13700 $D=4
M68 78 70 VSS VSS nch L=6e-08 W=1.5e-07 $X=48115 $Y=22800 $D=4
M69 VSS 85 83 VSS nch L=6e-08 W=2.6e-07 $X=48335 $Y=13665 $D=4
M70 32 87 VSS VSS nch L=6e-08 W=2.05e-07 $X=48570 $Y=10995 $D=4
M71 140 83 VSS VSS nch L=6e-08 W=1.5e-07 $X=48645 $Y=13700 $D=4
M72 VSS 87 32 VSS nch L=6e-08 W=2.05e-07 $X=48830 $Y=10995 $D=4
M73 85 89 140 VSS nch L=6e-08 W=1.5e-07 $X=48885 $Y=13700 $D=4
M74 87 clk VSS VSS nch L=6e-08 W=2.05e-07 $X=49090 $Y=10995 $D=4
M75 141 86 85 VSS nch L=6e-08 W=2.7e-07 $X=49160 $Y=13700 $D=4
M76 VSS 91 141 VSS nch L=6e-08 W=2.35e-07 $X=49390 $Y=13745 $D=4
M77 VSS 91 89 VSS nch L=6e-08 W=1.5e-07 $X=49855 $Y=13700 $D=4
M78 91 32 VSS VSS nch L=6e-08 W=1.5e-07 $X=50115 $Y=13700 $D=4
M79 142 82 70 VSS nch L=6e-08 W=3e-07 $X=50270 $Y=19300 $D=4
M80 143 93 142 VSS nch L=6e-08 W=3e-07 $X=50530 $Y=19300 $D=4
M81 144 94 143 VSS nch L=6e-08 W=3e-07 $X=50790 $Y=19300 $D=4
M82 VSS 88 144 VSS nch L=6e-08 W=3e-07 $X=51050 $Y=19300 $D=4
M83 VSS 95 81 VSS nch L=6e-08 W=2.8e-07 $X=51225 $Y=16500 $D=4
M84 VSS 97 95 VSS nch L=6e-08 W=1.9e-07 $X=51705 $Y=16465 $D=4
M85 96 95 VSS VSS nch L=6e-08 W=1.5e-07 $X=51955 $Y=16630 $D=4
M86 97 107 96 VSS nch L=6e-08 W=1.5e-07 $X=52295 $Y=16630 $D=4
M87 145 80 86 VSS nch L=6e-08 W=3e-07 $X=52450 $Y=11600 $D=4
M88 98 106 97 VSS nch L=6e-08 W=1.5e-07 $X=52600 $Y=16500 $D=4
M89 VSS 99 145 VSS nch L=6e-08 W=3e-07 $X=52710 $Y=11600 $D=4
M90 VSS 101 98 VSS nch L=6e-08 W=2.6e-07 $X=52935 $Y=16465 $D=4
M91 146 98 VSS VSS nch L=6e-08 W=1.5e-07 $X=53245 $Y=16500 $D=4
M92 101 106 146 VSS nch L=6e-08 W=1.5e-07 $X=53485 $Y=16500 $D=4
M93 147 102 101 VSS nch L=6e-08 W=2.7e-07 $X=53760 $Y=16500 $D=4
M94 VSS 107 147 VSS nch L=6e-08 W=2.35e-07 $X=53990 $Y=16545 $D=4
M95 VSS 107 106 VSS nch L=6e-08 W=1.5e-07 $X=54455 $Y=16500 $D=4
M96 107 32 VSS VSS nch L=6e-08 W=1.5e-07 $X=54715 $Y=16500 $D=4
M97 VDD 10 11 VDD pch L=6e-08 W=3.8e-07 $X=10250 $Y=10200 $D=103
M98 clk_out 11 VDD VDD pch L=6e-08 W=3.8e-07 $X=10630 $Y=10200 $D=103
M99 VDD 11 clk_out VDD pch L=6e-08 W=3.8e-07 $X=10890 $Y=10200 $D=103
M100 VDD 40 12 VDD pch L=6e-08 W=3.6e-07 $X=27030 $Y=13020 $D=103
M101 13 15 VDD VDD pch L=6e-08 W=3.25e-07 $X=27340 $Y=13020 $D=103
M102 VDD 17 15 VDD pch L=6e-08 W=1.9e-07 $X=27865 $Y=13155 $D=103
M103 40 15 VDD VDD pch L=6e-08 W=1.5e-07 $X=28115 $Y=13020 $D=103
M104 17 21 40 VDD pch L=6e-08 W=1.5e-07 $X=28405 $Y=13150 $D=103
M105 18 30 17 VDD pch L=6e-08 W=1.5e-07 $X=28665 $Y=13150 $D=103
M106 VDD 22 18 VDD pch L=6e-08 W=1.65e-07 $X=28985 $Y=13180 $D=103
M107 VDD 20 10 VDD pch L=6e-08 W=1.9e-07 $X=29015 $Y=10200 $D=103
M108 109 19 VDD VDD pch L=6e-08 W=1.9e-07 $X=29275 $Y=10200 $D=103
M109 110 18 VDD VDD pch L=6e-08 W=1.65e-07 $X=29365 $Y=13180 $D=103
M110 20 27 109 VDD pch L=6e-08 W=1.6e-07 $X=29500 $Y=10200 $D=103
M111 22 30 110 VDD pch L=6e-08 W=1.5e-07 $X=29640 $Y=13100 $D=103
M112 111 26 20 VDD pch L=6e-08 W=1.6e-07 $X=29775 $Y=10200 $D=103
M113 39 21 22 VDD pch L=6e-08 W=1.65e-07 $X=29920 $Y=13180 $D=103
M114 VDD clk 111 VDD pch L=6e-08 W=1.8e-07 $X=30035 $Y=10400 $D=103
M115 VDD 37 25 VDD pch L=6e-08 W=3.6e-07 $X=30230 $Y=24220 $D=103
M116 27 26 VDD VDD pch L=6e-08 W=1.9e-07 $X=30315 $Y=10390 $D=103
M117 VDD 30 21 VDD pch L=6e-08 W=1.9e-07 $X=30410 $Y=13155 $D=103
M118 31 36 VDD VDD pch L=6e-08 W=3.25e-07 $X=30540 $Y=24220 $D=103
M119 30 32 VDD VDD pch L=6e-08 W=1.9e-07 $X=30650 $Y=13155 $D=103
M120 VDD 38 36 VDD pch L=6e-08 W=2e-07 $X=31080 $Y=24345 $D=103
M121 VDD 28 39 VDD pch L=6e-08 W=1.5e-07 $X=31230 $Y=13200 $D=103
M122 37 36 VDD VDD pch L=6e-08 W=1.9e-07 $X=31330 $Y=24310 $D=103
M123 38 46 37 VDD pch L=6e-08 W=1.5e-07 $X=31620 $Y=24350 $D=103
M124 112 12 VDD VDD pch L=6e-08 W=3.5e-07 $X=31640 $Y=13000 $D=103
M125 39 43 112 VDD pch L=6e-08 W=3.5e-07 $X=31840 $Y=13000 $D=103
M126 42 48 38 VDD pch L=6e-08 W=1.5e-07 $X=31920 $Y=24350 $D=103
M127 113 40 39 VDD pch L=6e-08 W=1.7e-07 $X=32180 $Y=13020 $D=103
M128 VDD 44 42 VDD pch L=6e-08 W=3.25e-07 $X=32265 $Y=24220 $D=103
M129 VDD 47 113 VDD pch L=6e-08 W=1.7e-07 $X=32405 $Y=13020 $D=103
M130 114 42 VDD VDD pch L=6e-08 W=1.5e-07 $X=32585 $Y=24350 $D=103
M131 43 47 VDD VDD pch L=6e-08 W=1.5e-07 $X=32715 $Y=13155 $D=103
M132 44 48 114 VDD pch L=6e-08 W=1.5e-07 $X=32810 $Y=24350 $D=103
M133 45 46 44 VDD pch L=6e-08 W=1.95e-07 $X=33195 $Y=24220 $D=103
M134 VDD 28 45 VDD pch L=6e-08 W=3.6e-07 $X=33540 $Y=24220 $D=103
M135 45 25 VDD VDD pch L=6e-08 W=1.9e-07 $X=33780 $Y=24390 $D=103
M136 VDD 48 46 VDD pch L=6e-08 W=1.9e-07 $X=34270 $Y=24390 $D=103
M137 48 32 VDD VDD pch L=6e-08 W=1.9e-07 $X=34515 $Y=24390 $D=103
M138 VDD 50 52 VDD pch L=6e-08 W=2.7e-07 $X=38415 $Y=17820 $D=103
M139 115 49 VDD VDD pch L=6e-08 W=1.8e-07 $X=38700 $Y=17820 $D=103
M140 55 50 115 VDD pch L=6e-08 W=2.2e-07 $X=38955 $Y=17980 $D=103
M141 56 34 VDD VDD pch L=6e-08 W=1.9e-07 $X=39235 $Y=21420 $D=103
M142 116 52 55 VDD pch L=6e-08 W=2.1e-07 $X=39250 $Y=17820 $D=103
M143 VDD 53 116 VDD pch L=6e-08 W=2.1e-07 $X=39455 $Y=17820 $D=103
M144 VDD 51 56 VDD pch L=6e-08 W=1.9e-07 $X=39475 $Y=21550 $D=103
M145 60 55 VDD VDD pch L=6e-08 W=2.95e-07 $X=39725 $Y=17905 $D=103
M146 117 54 VDD VDD pch L=6e-08 W=1.9e-07 $X=39735 $Y=21550 $D=103
M147 56 60 117 VDD pch L=6e-08 W=1.9e-07 $X=39925 $Y=21550 $D=103
M148 VDD 74 68 VDD pch L=6e-08 W=3.6e-07 $X=46225 $Y=13020 $D=103
M149 69 72 VDD VDD pch L=6e-08 W=3.25e-07 $X=46540 $Y=13020 $D=103
M150 118 68 76 VDD pch L=6e-08 W=3.8e-07 $X=46830 $Y=17820 $D=103
M151 VDD 75 63 VDD pch L=6e-08 W=3.8e-07 $X=47015 $Y=15020 $D=103
M152 VDD 79 72 VDD pch L=6e-08 W=1.9e-07 $X=47080 $Y=13155 $D=103
M153 119 66 118 VDD pch L=6e-08 W=3.8e-07 $X=47080 $Y=17820 $D=103
M154 75 69 VDD VDD pch L=6e-08 W=1.85e-07 $X=47285 $Y=15020 $D=103
M155 VDD 26 71 VDD pch L=6e-08 W=1.9e-07 $X=47285 $Y=23610 $D=103
M156 74 72 VDD VDD pch L=6e-08 W=1.5e-07 $X=47330 $Y=13150 $D=103
M157 120 53 119 VDD pch L=6e-08 W=3.8e-07 $X=47330 $Y=17820 $D=103
M158 VDD 77 75 VDD pch L=6e-08 W=1.85e-07 $X=47545 $Y=15020 $D=103
M159 VDD 65 120 VDD pch L=6e-08 W=3.8e-07 $X=47580 $Y=17820 $D=103
M160 121 71 VDD VDD pch L=6e-08 W=3.8e-07 $X=47595 $Y=23420 $D=103
M161 79 89 74 VDD pch L=6e-08 W=1.5e-07 $X=47620 $Y=13150 $D=103
M162 122 77 121 VDD pch L=6e-08 W=3.8e-07 $X=47855 $Y=23420 $D=103
M163 26 76 VDD VDD pch L=6e-08 W=3.8e-07 $X=47860 $Y=17820 $D=103
M164 83 91 79 VDD pch L=6e-08 W=1.5e-07 $X=48000 $Y=13150 $D=103
M165 78 70 122 VDD pch L=6e-08 W=3.8e-07 $X=48115 $Y=23420 $D=103
M166 VDD 85 83 VDD pch L=6e-08 W=3.25e-07 $X=48335 $Y=13020 $D=103
M167 32 87 VDD VDD pch L=6e-08 W=3.8e-07 $X=48570 $Y=10200 $D=103
M168 123 83 VDD VDD pch L=6e-08 W=1.5e-07 $X=48645 $Y=13150 $D=103
M169 VDD 87 32 VDD pch L=6e-08 W=3.8e-07 $X=48830 $Y=10200 $D=103
M170 85 91 123 VDD pch L=6e-08 W=1.5e-07 $X=48885 $Y=13150 $D=103
M171 87 clk VDD VDD pch L=6e-08 W=3.8e-07 $X=49115 $Y=10200 $D=103
M172 124 86 85 VDD pch L=6e-08 W=3.5e-07 $X=49160 $Y=13020 $D=103
M173 VDD 89 124 VDD pch L=6e-08 W=2.75e-07 $X=49395 $Y=13020 $D=103
M174 VDD 91 89 VDD pch L=6e-08 W=1.9e-07 $X=49870 $Y=13190 $D=103
M175 91 32 VDD VDD pch L=6e-08 W=1.9e-07 $X=50115 $Y=13190 $D=103
M176 70 82 VDD VDD pch L=6e-08 W=3.8e-07 $X=50270 $Y=18600 $D=103
M177 VDD 93 70 VDD pch L=6e-08 W=3.8e-07 $X=50530 $Y=18600 $D=103
M178 70 94 VDD VDD pch L=6e-08 W=3.8e-07 $X=50790 $Y=18600 $D=103
M179 VDD 88 70 VDD pch L=6e-08 W=3.8e-07 $X=51050 $Y=18600 $D=103
M180 VDD 95 81 VDD pch L=6e-08 W=3.25e-07 $X=51220 $Y=15820 $D=103
M181 VDD 97 95 VDD pch L=6e-08 W=1.9e-07 $X=51680 $Y=15955 $D=103
M182 96 95 VDD VDD pch L=6e-08 W=1.5e-07 $X=51930 $Y=15950 $D=103
M183 97 106 96 VDD pch L=6e-08 W=1.5e-07 $X=52220 $Y=15950 $D=103
M184 86 80 VDD VDD pch L=6e-08 W=3.8e-07 $X=52450 $Y=12220 $D=103
M185 98 107 97 VDD pch L=6e-08 W=1.5e-07 $X=52600 $Y=15950 $D=103
M186 VDD 99 86 VDD pch L=6e-08 W=3.8e-07 $X=52710 $Y=12220 $D=103
M187 VDD 101 98 VDD pch L=6e-08 W=3.25e-07 $X=52935 $Y=15820 $D=103
M188 125 98 VDD VDD pch L=6e-08 W=1.5e-07 $X=53245 $Y=15950 $D=103
M189 101 107 125 VDD pch L=6e-08 W=1.5e-07 $X=53485 $Y=15950 $D=103
M190 126 102 101 VDD pch L=6e-08 W=3.5e-07 $X=53760 $Y=15820 $D=103
M191 VDD 106 126 VDD pch L=6e-08 W=2.75e-07 $X=53995 $Y=15820 $D=103
M192 VDD 107 106 VDD pch L=6e-08 W=1.9e-07 $X=54470 $Y=15990 $D=103
M193 107 32 VDD VDD pch L=6e-08 W=1.9e-07 $X=54715 $Y=15990 $D=103
X237 VSS VDD ICV_11 $T=49800 11400 1 0 $X=49565 $Y=9765
X238 VSS VDD DCAP4BWP7T $T=30000 22600 1 0 $X=29765 $Y=20965
X239 VSS VDD DCAP4BWP7T $T=35600 19800 0 0 $X=35365 $Y=19695
X240 VSS VDD DCAP4BWP7T $T=37600 19800 0 0 $X=37365 $Y=19695
X241 VSS VDD DCAP4BWP7T $T=37600 22600 1 0 $X=37365 $Y=20965
X242 VSS VDD DCAP4BWP7T $T=40400 19800 1 0 $X=40165 $Y=18165
X243 VSS VDD DCAP4BWP7T $T=43800 14200 1 0 $X=43565 $Y=12565
X244 VSS VDD DCAP4BWP7T $T=43800 17000 1 0 $X=43565 $Y=15365
X245 VSS VDD DCAP4BWP7T $T=47800 14200 0 0 $X=47565 $Y=14095
X246 VSS VDD DCAP4BWP7T $T=48200 17000 0 0 $X=47965 $Y=16895
X247 VSS VDD DCAP4BWP7T $T=51400 14200 0 0 $X=51165 $Y=14095
X248 VSS VDD DCAP4BWP7T $T=55600 11400 1 0 $X=55365 $Y=9765
X249 VSS VDD DCAP4BWP7T $T=55600 14200 1 0 $X=55365 $Y=12565
X250 VSS VDD DCAP4BWP7T $T=55600 17000 1 0 $X=55365 $Y=15365
X251 VSS VDD DCAP4BWP7T $T=55600 22600 1 0 $X=55365 $Y=20965
X252 VSS VDD DCAP4BWP7T $T=55600 25400 0 0 $X=55365 $Y=25295
X253 VSS VDD DCAP4BWP7T $T=58800 14200 0 0 $X=58565 $Y=14095
X262 VSS VDD ICV_9 $T=44200 22600 1 0 $X=43965 $Y=20965
X263 VSS VDD ICV_9 $T=54200 25400 0 0 $X=53965 $Y=25295
X264 VDD VSS DCAP32BWP7T $T=48400 22600 0 0 $X=48165 $Y=22495
X265 VDD VSS DCAP8BWP7T $T=13400 11400 1 0 $X=13165 $Y=9765
X266 VDD VSS DCAP8BWP7T $T=26600 11400 1 0 $X=26365 $Y=9765
X267 VDD VSS DCAP8BWP7T $T=32000 19800 0 0 $X=31765 $Y=19695
X268 VDD VSS DCAP8BWP7T $T=36000 22600 1 0 $X=35765 $Y=20965
X269 VDD VSS DCAP8BWP7T $T=38400 19800 0 0 $X=38165 $Y=19695
X270 VDD VSS DCAP8BWP7T $T=52200 14200 0 0 $X=51965 $Y=14095
X271 VDD VSS DCAP8BWP7T $T=53400 11400 1 0 $X=53165 $Y=9765
X272 VDD VSS DCAP8BWP7T $T=56200 22600 0 0 $X=55965 $Y=22495
X273 VSS VDD ICV_1 $T=33600 14200 0 0 $X=33365 $Y=14095
X274 VSS VDD ICV_1 $T=33600 19800 0 0 $X=33365 $Y=19695
X275 VSS VDD ICV_1 $T=34000 11400 1 0 $X=33765 $Y=9765
X276 VSS VDD ICV_1 $T=35600 14200 0 0 $X=35365 $Y=14095
X277 VSS VDD ICV_1 $T=37400 19800 1 0 $X=37165 $Y=18165
X278 VSS VDD ICV_1 $T=45600 17000 1 0 $X=45365 $Y=15365
X279 VSS VDD ICV_1 $T=46000 22600 0 0 $X=45765 $Y=22495
X280 VSS VDD ICV_1 $T=53800 25400 1 0 $X=53565 $Y=23765
X281 VSS VDD ICV_1 $T=58600 22600 0 0 $X=58365 $Y=22495
X282 VDD VSS ICV_12 $T=16000 11400 1 0 $X=15765 $Y=9765
X283 VDD VSS ICV_12 $T=45800 28200 1 0 $X=45565 $Y=26565
X284 VDD VSS ICV_12 $T=45800 28200 0 0 $X=45565 $Y=28095
X285 VDD VSS ICV_12 $T=45800 31000 1 0 $X=45565 $Y=29365
X286 VDD VSS ICV_12 $T=45800 31000 0 0 $X=45565 $Y=30895
X287 VDD VSS ICV_12 $T=45800 33800 1 0 $X=45565 $Y=32165
X288 VSS VDD ICV_19 $T=10000 11400 0 0 $X=9765 $Y=11295
X289 VSS VDD ICV_19 $T=10000 14200 0 0 $X=9765 $Y=14095
X290 VSS VDD ICV_19 $T=10000 17000 0 0 $X=9765 $Y=16895
X291 VSS VDD ICV_19 $T=10000 19800 0 0 $X=9765 $Y=19695
X292 VSS VDD ICV_19 $T=10000 22600 0 0 $X=9765 $Y=22495
X293 VSS VDD ICV_19 $T=10000 25400 0 0 $X=9765 $Y=25295
X294 VSS VDD ICV_19 $T=10000 28200 0 0 $X=9765 $Y=28095
X295 VSS VDD ICV_19 $T=10000 31000 0 0 $X=9765 $Y=30895
X296 VSS VDD ICV_4 $T=11600 11400 1 0 $X=11365 $Y=9765
X297 VSS VDD ICV_4 $T=26600 17000 0 0 $X=26365 $Y=16895
X298 VSS VDD ICV_4 $T=36000 11400 1 0 $X=35765 $Y=9765
X299 VSS VDD ICV_4 $T=41400 19800 0 0 $X=41165 $Y=19695
X300 VSS VDD ICV_4 $T=56200 11400 0 0 $X=55965 $Y=11295
X301 VSS VDD ICV_13 $T=25000 11400 1 0 $X=24765 $Y=9765
X302 VSS VDD ICV_13 $T=25000 14200 1 0 $X=24765 $Y=12565
X303 VSS VDD ICV_13 $T=25000 17000 1 0 $X=24765 $Y=15365
X304 VSS VDD ICV_13 $T=25000 17000 0 0 $X=24765 $Y=16895
X305 VSS VDD ICV_13 $T=25000 19800 1 0 $X=24765 $Y=18165
X306 VSS VDD ICV_13 $T=25000 19800 0 0 $X=24765 $Y=19695
X307 VSS VDD ICV_13 $T=25000 22600 1 0 $X=24765 $Y=20965
X308 VSS VDD ICV_13 $T=25000 25400 1 0 $X=24765 $Y=23765
X309 VSS VDD ICV_13 $T=45000 11400 1 0 $X=44765 $Y=9765
X310 VSS VDD ICV_10 $T=25600 14200 0 0 $X=25365 $Y=14095
X311 VSS VDD ICV_10 $T=31800 14200 0 0 $X=31565 $Y=14095
X312 VSS VDD ICV_10 $T=31800 19800 1 0 $X=31565 $Y=18165
X313 VSS VDD ICV_10 $T=41000 14200 0 0 $X=40765 $Y=14095
X314 VSS VDD ICV_10 $T=45600 22600 1 0 $X=45365 $Y=20965
X315 VSS VDD ICV_10 $T=52000 25400 1 0 $X=51765 $Y=23765
X318 VDD VSS ICV_15 $T=36200 25400 1 0 $X=35965 $Y=23765
X319 VSS VDD ICV_16 $T=25000 11400 0 0 $X=24765 $Y=11295
X320 VSS VDD ICV_16 $T=25000 22600 0 0 $X=24765 $Y=22495
X321 VSS VDD ICV_16 $T=25000 25400 0 0 $X=24765 $Y=25295
X322 VSS VDD ICV_16 $T=25000 28200 1 0 $X=24765 $Y=26565
X323 VSS VDD ICV_16 $T=25000 28200 0 0 $X=24765 $Y=28095
X324 VSS VDD ICV_16 $T=25000 31000 1 0 $X=24765 $Y=29365
X325 VSS VDD ICV_16 $T=25000 31000 0 0 $X=24765 $Y=30895
X326 VSS VDD ICV_16 $T=25000 33800 1 0 $X=24765 $Y=32165
X345 VSS VDD ICV_2 $T=26600 22600 1 0 $X=26365 $Y=20965
X346 VSS VDD ICV_2 $T=26600 25400 1 0 $X=26365 $Y=23765
X347 VSS VDD ICV_2 $T=30600 11400 1 0 $X=30365 $Y=9765
X348 32 16 28 VDD VSS 14 DFKCNQD1BWP7T $T=31800 14200 1 180 $X=27165 $Y=14095
X349 32 57 28 VDD VSS 50 DFKCNQD1BWP7T $T=41000 14200 1 180 $X=36365 $Y=14095
X350 32 100 99 VDD VSS 84 DFKCNQD1BWP7T $T=54600 22600 0 180 $X=49965 $Y=20965
X351 32 103 99 VDD VSS 90 DFKCNQD1BWP7T $T=54800 19800 1 180 $X=50165 $Y=19695
X352 32 104 99 VDD VSS 92 DFKCNQD1BWP7T $T=55000 14200 0 180 $X=50365 $Y=12565
X376 35 31 14 VSS VDD 16 HA1D0BWP7T $T=31400 17000 1 180 $X=28165 $Y=16895
X377 47 50 35 VSS VDD 57 HA1D0BWP7T $T=37200 17000 1 0 $X=36965 $Y=15365
X378 67 65 62 VSS VDD 24 HA1D0BWP7T $T=44200 19800 0 180 $X=40965 $Y=18165
X379 62 66 63 VSS VDD 29 HA1D0BWP7T $T=44400 17000 1 180 $X=41165 $Y=16895
X380 35 29 24 23 12 VDD VSS OAI31D1BWP7T $T=31000 19800 0 180 $X=29365 $Y=18165
X381 div_sel[2] 100 div_sel[1] 105 108 VDD VSS OAI31D1BWP7T $T=57400 14200 0 0 $X=57165 $Y=14095
X382 24 34 33 23 VDD VSS AOI21D0BWP7T $T=31400 19800 1 180 $X=30165 $Y=19695
X383 54 59 58 56 VDD VSS AOI21D0BWP7T $T=41000 19800 1 180 $X=39765 $Y=19695
X384 31 14 33 29 VSS VDD MUX2ND0BWP7T $T=30800 22600 1 0 $X=30565 $Y=20965
X385 69 73 80 81 VSS VDD MUX2ND0BWP7T $T=46600 11400 1 0 $X=46365 $Y=9765
X401 24 VSS 49 14 VDD IND2D1BWP7T $T=37400 19800 0 180 $X=36165 $Y=18165
X402 59 VSS 64 26 VDD IND2D1BWP7T $T=43200 19800 0 0 $X=42965 $Y=19695
X403 49 25 VSS 51 29 VDD IOA21D0BWP7T $T=36400 19800 0 0 $X=36165 $Y=19695
X404 59 70 VSS 73 26 VDD IOA21D0BWP7T $T=46400 19800 0 0 $X=46165 $Y=19695
X405 64 61 rst_n 32 VSS VDD 19 EDFKCNQD1BWP7T $T=43600 11400 0 180 $X=37565 $Y=9765
X406 73 84 rst_n 32 VSS VDD 53 EDFKCNQD1BWP7T $T=51800 25400 1 180 $X=45765 $Y=25295
X407 64 78 rst_n 32 VSS VDD 77 EDFKCNQD1BWP7T $T=46200 25400 1 0 $X=45965 $Y=23765
X408 73 92 rst_n 32 VSS VDD 66 EDFKCNQD1BWP7T $T=52200 11400 1 180 $X=46165 $Y=11295
X409 73 90 rst_n 32 VSS VDD 65 EDFKCNQD1BWP7T $T=49000 17000 0 0 $X=48765 $Y=16895
X410 49 50 VDD VSS 58 XOR2D1BWP7T $T=38400 19800 1 0 $X=38165 $Y=18165
X411 67 53 VDD VSS 54 XOR2D1BWP7T $T=44200 22600 0 180 $X=41965 $Y=20965
X412 26 VDD 61 19 VSS INR2XD0BWP7T $T=43800 14200 0 180 $X=42565 $Y=12565
X413 rst_n VDD 28 64 VSS INR2XD0BWP7T $T=42800 14200 0 0 $X=42565 $Y=14095
X414 rst_n VDD 108 div_sel[0] VSS INR2XD0BWP7T $T=58000 11400 0 0 $X=57765 $Y=11295
X415 69 81 VDD VSS 82 XNR2D1BWP7T $T=46600 17000 1 0 $X=46365 $Y=15365
X416 53 84 VDD VSS 88 XNR2D1BWP7T $T=47400 22600 1 0 $X=47165 $Y=20965
X417 66 92 VDD VSS 93 XNR2D1BWP7T $T=49000 14200 0 0 $X=48765 $Y=14095
X418 65 90 VDD VSS 94 XNR2D1BWP7T $T=54800 19800 0 180 $X=52565 $Y=18165
X419 rst_n VSS VDD 99 BUFFD1BWP7T $T=53400 25400 0 0 $X=53165 $Y=25295
X420 105 VSS VDD 102 BUFFD1BWP7T $T=53800 14200 0 0 $X=53565 $Y=14095
X421 div_sel[1] VSS VDD 104 BUFFD1BWP7T $T=54000 11400 0 0 $X=53765 $Y=11295
X422 div_sel[2] VSS VDD 103 BUFFD1BWP7T $T=55600 19800 0 0 $X=55365 $Y=19695
X423 div_sel[3] VSS VDD 100 BUFFD1BWP7T $T=57800 22600 0 0 $X=57565 $Y=22495
X424 VSS VDD ICV_3 $T=56400 11400 1 0 $X=56165 $Y=9765
X425 VSS VDD ICV_3 $T=56400 17000 1 0 $X=56165 $Y=15365
X426 VSS VDD ICV_3 $T=56400 19800 0 0 $X=56165 $Y=19695
X427 VSS VDD ICV_3 $T=56400 22600 1 0 $X=56165 $Y=20965
X428 VSS VDD ICV_3 $T=56400 25400 0 0 $X=56165 $Y=25295
X429 VSS VDD ICV_7 $T=54800 17000 0 0 $X=54565 $Y=16895
X430 VSS VDD ICV_7 $T=54800 19800 1 0 $X=54565 $Y=18165
X431 VSS VDD ICV_7 $T=54800 25400 1 0 $X=54565 $Y=23765
X432 VSS VDD ICV_7 $T=54800 28200 1 0 $X=54565 $Y=26565
X433 VSS VDD ICV_7 $T=54800 28200 0 0 $X=54565 $Y=28095
X434 VSS VDD ICV_7 $T=54800 31000 1 0 $X=54565 $Y=29365
X435 VSS VDD ICV_7 $T=54800 31000 0 0 $X=54565 $Y=30895
X436 VSS VDD ICV_7 $T=54800 33800 1 0 $X=54565 $Y=32165
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410915 1
** N=1 EP=1 IP=0 FDC=5
M0 1 1 1 1 nch L=2e-07 W=2e-06 $X=0 $Y=0 $D=4
M1 1 1 1 1 nch L=2e-07 W=2e-06 $X=400 $Y=0 $D=4
M2 1 1 1 1 nch L=2e-07 W=2e-06 $X=800 $Y=0 $D=4
M3 1 1 1 1 nch L=2e-07 W=2e-06 $X=1200 $Y=0 $D=4
M4 1 1 1 1 nch L=2e-07 W=2e-06 $X=1600 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410912 1 2 3 4
** N=4 EP=4 IP=0 FDC=5
M0 2 3 1 4 nch L=2e-07 W=2e-06 $X=0 $Y=0 $D=4
M1 1 3 2 4 nch L=2e-07 W=2e-06 $X=400 $Y=0 $D=4
M2 2 3 1 4 nch L=2e-07 W=2e-06 $X=800 $Y=0 $D=4
M3 1 3 2 4 nch L=2e-07 W=2e-06 $X=1200 $Y=0 $D=4
M4 2 3 1 4 nch L=2e-07 W=2e-06 $X=1600 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT pch_CDNS_7649669410911 1
** N=2 EP=1 IP=0 FDC=2
M0 1 1 1 1 pch L=1.5e-07 W=4.5e-06 $X=0 $Y=0 $D=103
M1 1 1 1 1 pch L=1.5e-07 W=4.5e-06 $X=350 $Y=0 $D=103
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410914 1
** N=1 EP=1 IP=0 FDC=2
M0 1 1 1 1 nch L=1.5e-07 W=2e-06 $X=0 $Y=0 $D=4
M1 1 1 1 1 nch L=1.5e-07 W=2e-06 $X=350 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT pch_CDNS_764966941092 1 2 3 5
** N=5 EP=4 IP=0 FDC=2
M0 2 3 1 5 pch L=1.5e-07 W=4.5e-06 $X=0 $Y=0 $D=103
M1 1 3 2 5 pch L=1.5e-07 W=4.5e-06 $X=350 $Y=0 $D=103
.ENDS
***************************************
.SUBCKT nch_CDNS_764966941093 1 2 3 4
** N=4 EP=4 IP=0 FDC=2
M0 2 3 1 4 nch L=1.5e-07 W=2e-06 $X=0 $Y=0 $D=4
M1 1 3 2 4 nch L=1.5e-07 W=2e-06 $X=350 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT pch_lvt_CDNS_764966941098 1
** N=2 EP=1 IP=0 FDC=10
M0 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=0 $Y=0 $D=121
M1 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=260 $Y=0 $D=121
M2 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=520 $Y=0 $D=121
M3 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=780 $Y=0 $D=121
M4 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=1040 $Y=0 $D=121
M5 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=1300 $Y=0 $D=121
M6 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=1560 $Y=0 $D=121
M7 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=1820 $Y=0 $D=121
M8 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=2080 $Y=0 $D=121
M9 1 1 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=2340 $Y=0 $D=121
.ENDS
***************************************
.SUBCKT nch_lvt_CDNS_764966941099 1
** N=1 EP=1 IP=0 FDC=10
M0 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=0 $Y=0 $D=45
M1 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=260 $Y=0 $D=45
M2 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=520 $Y=0 $D=45
M3 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=780 $Y=0 $D=45
M4 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=1040 $Y=0 $D=45
M5 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=1300 $Y=0 $D=45
M6 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=1560 $Y=0 $D=45
M7 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=1820 $Y=0 $D=45
M8 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=2080 $Y=0 $D=45
M9 1 1 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=2340 $Y=0 $D=45
.ENDS
***************************************
.SUBCKT pch_lvt_CDNS_7649669410913 1 2 3
** N=4 EP=3 IP=0 FDC=10
M0 2 3 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=0 $Y=0 $D=121
M1 1 3 2 1 pch_lvt L=6e-08 W=4.56e-06 $X=260 $Y=0 $D=121
M2 2 3 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=520 $Y=0 $D=121
M3 1 3 2 1 pch_lvt L=6e-08 W=4.56e-06 $X=780 $Y=0 $D=121
M4 2 3 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=1040 $Y=0 $D=121
M5 1 3 2 1 pch_lvt L=6e-08 W=4.56e-06 $X=1300 $Y=0 $D=121
M6 2 3 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=1560 $Y=0 $D=121
M7 1 3 2 1 pch_lvt L=6e-08 W=4.56e-06 $X=1820 $Y=0 $D=121
M8 2 3 1 1 pch_lvt L=6e-08 W=4.56e-06 $X=2080 $Y=0 $D=121
M9 1 3 2 1 pch_lvt L=6e-08 W=4.56e-06 $X=2340 $Y=0 $D=121
.ENDS
***************************************
.SUBCKT nch_lvt_CDNS_7649669410910 1 2 3
** N=3 EP=3 IP=0 FDC=10
M0 2 3 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=0 $Y=0 $D=45
M1 1 3 2 1 nch_lvt L=6e-08 W=3.6e-06 $X=260 $Y=0 $D=45
M2 2 3 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=520 $Y=0 $D=45
M3 1 3 2 1 nch_lvt L=6e-08 W=3.6e-06 $X=780 $Y=0 $D=45
M4 2 3 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=1040 $Y=0 $D=45
M5 1 3 2 1 nch_lvt L=6e-08 W=3.6e-06 $X=1300 $Y=0 $D=45
M6 2 3 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=1560 $Y=0 $D=45
M7 1 3 2 1 nch_lvt L=6e-08 W=3.6e-06 $X=1820 $Y=0 $D=45
M8 2 3 1 1 nch_lvt L=6e-08 W=3.6e-06 $X=2080 $Y=0 $D=45
M9 1 3 2 1 nch_lvt L=6e-08 W=3.6e-06 $X=2340 $Y=0 $D=45
.ENDS
***************************************
.SUBCKT Ring_VCO vctrl VDD VSS f_out
** N=23 EP=4 IP=236 FDC=516
M0 VSS 7 7 VSS nch L=1e-06 W=2e-06 $X=39000 $Y=-11705 $D=4
M1 6 6 VDD VDD pch L=3e-07 W=4.5e-06 $X=35950 $Y=-4605 $D=103
M2 VDD 6 7 VDD pch L=1e-06 W=4.5e-06 $X=39000 $Y=-4605 $D=103
X3 5 VSS rpodwo l=2e-05 w=4.5e-07 $X=48795 $Y=-34790 $D=476
X4 VSS nch_CDNS_7649669410915 $T=23230 -34130 0 0 $X=22925 $Y=-34470
X5 VSS nch_CDNS_7649669410915 $T=23230 -29050 0 0 $X=22925 $Y=-29390
X6 VSS nch_CDNS_7649669410915 $T=23230 -23970 0 0 $X=22925 $Y=-24310
X7 VSS nch_CDNS_7649669410915 $T=23230 -18890 0 0 $X=22925 $Y=-19230
X8 VSS nch_CDNS_7649669410915 $T=28220 -34130 0 0 $X=27915 $Y=-34470
X9 VSS nch_CDNS_7649669410915 $T=28220 -18890 0 0 $X=27915 $Y=-19230
X10 VSS nch_CDNS_7649669410915 $T=33210 -34130 0 0 $X=32905 $Y=-34470
X11 VSS nch_CDNS_7649669410915 $T=33210 -18890 0 0 $X=32905 $Y=-19230
X12 VSS nch_CDNS_7649669410915 $T=38200 -34130 0 0 $X=37895 $Y=-34470
X13 VSS nch_CDNS_7649669410915 $T=38200 -29050 0 0 $X=37895 $Y=-29390
X14 VSS nch_CDNS_7649669410915 $T=38200 -23970 0 0 $X=37895 $Y=-24310
X15 VSS nch_CDNS_7649669410915 $T=38200 -18890 0 0 $X=37895 $Y=-19230
X16 5 6 vctrl VSS nch_CDNS_7649669410912 $T=28220 -29050 0 0 $X=27915 $Y=-29390
X17 5 6 vctrl VSS nch_CDNS_7649669410912 $T=28220 -23970 0 0 $X=27915 $Y=-24310
X18 5 6 vctrl VSS nch_CDNS_7649669410912 $T=33210 -29050 0 0 $X=32905 $Y=-29390
X19 5 6 vctrl VSS nch_CDNS_7649669410912 $T=33210 -23970 0 0 $X=32905 $Y=-24310
X20 VDD pch_CDNS_7649669410911 $T=48220 -4605 0 0 $X=47825 $Y=-4945
X21 VDD pch_CDNS_7649669410911 $T=48220 2575 0 0 $X=47825 $Y=2235
X22 VDD pch_CDNS_7649669410911 $T=48220 9755 0 0 $X=47825 $Y=9415
X23 VDD pch_CDNS_7649669410911 $T=48220 16935 0 0 $X=47825 $Y=16595
X24 VDD pch_CDNS_7649669410911 $T=51510 -4605 0 0 $X=51115 $Y=-4945
X25 VDD pch_CDNS_7649669410911 $T=51510 16935 0 0 $X=51115 $Y=16595
X26 VDD pch_CDNS_7649669410911 $T=54800 -4605 0 0 $X=54405 $Y=-4945
X27 VDD pch_CDNS_7649669410911 $T=54800 16935 0 0 $X=54405 $Y=16595
X28 VDD pch_CDNS_7649669410911 $T=58090 -4605 0 0 $X=57695 $Y=-4945
X29 VDD pch_CDNS_7649669410911 $T=58090 16935 0 0 $X=57695 $Y=16595
X30 VDD pch_CDNS_7649669410911 $T=61380 -4605 0 0 $X=60985 $Y=-4945
X31 VDD pch_CDNS_7649669410911 $T=61380 16935 0 0 $X=60985 $Y=16595
X32 VDD pch_CDNS_7649669410911 $T=64670 -4605 0 0 $X=64275 $Y=-4945
X33 VDD pch_CDNS_7649669410911 $T=64670 16935 0 0 $X=64275 $Y=16595
X34 VDD pch_CDNS_7649669410911 $T=67960 -4605 0 0 $X=67565 $Y=-4945
X35 VDD pch_CDNS_7649669410911 $T=67960 2575 0 0 $X=67565 $Y=2235
X36 VDD pch_CDNS_7649669410911 $T=67960 9755 0 0 $X=67565 $Y=9415
X37 VDD pch_CDNS_7649669410911 $T=67960 16935 0 0 $X=67565 $Y=16595
X38 VSS nch_CDNS_7649669410914 $T=48390 -27340 0 0 $X=48085 $Y=-27680
X39 VSS nch_CDNS_7649669410914 $T=48390 -22660 0 0 $X=48085 $Y=-23000
X40 VSS nch_CDNS_7649669410914 $T=48390 -17980 0 0 $X=48085 $Y=-18320
X41 VSS nch_CDNS_7649669410914 $T=48390 -13300 0 0 $X=48085 $Y=-13640
X42 VSS nch_CDNS_7649669410914 $T=51680 -27340 0 0 $X=51375 $Y=-27680
X43 VSS nch_CDNS_7649669410914 $T=51680 -13300 0 0 $X=51375 $Y=-13640
X44 VSS nch_CDNS_7649669410914 $T=54970 -27340 0 0 $X=54665 $Y=-27680
X45 VSS nch_CDNS_7649669410914 $T=54970 -13300 0 0 $X=54665 $Y=-13640
X46 VSS nch_CDNS_7649669410914 $T=58260 -27340 0 0 $X=57955 $Y=-27680
X47 VSS nch_CDNS_7649669410914 $T=58260 -13300 0 0 $X=57955 $Y=-13640
X48 VSS nch_CDNS_7649669410914 $T=61550 -27340 0 0 $X=61245 $Y=-27680
X49 VSS nch_CDNS_7649669410914 $T=61550 -13300 0 0 $X=61245 $Y=-13640
X50 VSS nch_CDNS_7649669410914 $T=64840 -27340 0 0 $X=64535 $Y=-27680
X51 VSS nch_CDNS_7649669410914 $T=64840 -13300 0 0 $X=64535 $Y=-13640
X52 VSS nch_CDNS_7649669410914 $T=68130 -27340 0 0 $X=67825 $Y=-27680
X53 VSS nch_CDNS_7649669410914 $T=68130 -22660 0 0 $X=67825 $Y=-23000
X54 VSS nch_CDNS_7649669410914 $T=68130 -17980 0 0 $X=67825 $Y=-18320
X55 VSS nch_CDNS_7649669410914 $T=68130 -13300 0 0 $X=67825 $Y=-13640
X56 10 8 9 VDD pch_CDNS_764966941092 $T=51510 2575 0 0 $X=51115 $Y=2235
X57 VDD 10 6 VDD pch_CDNS_764966941092 $T=51510 9755 0 0 $X=51115 $Y=9415
X58 13 12 8 VDD pch_CDNS_764966941092 $T=54800 2575 0 0 $X=54405 $Y=2235
X59 VDD 13 6 VDD pch_CDNS_764966941092 $T=54800 9755 0 0 $X=54405 $Y=9415
X60 16 15 12 VDD pch_CDNS_764966941092 $T=58090 2575 0 0 $X=57695 $Y=2235
X61 VDD 16 6 VDD pch_CDNS_764966941092 $T=58090 9755 0 0 $X=57695 $Y=9415
X62 19 18 15 VDD pch_CDNS_764966941092 $T=61380 2575 0 0 $X=60985 $Y=2235
X63 VDD 19 6 VDD pch_CDNS_764966941092 $T=61380 9755 0 0 $X=60985 $Y=9415
X64 21 9 18 VDD pch_CDNS_764966941092 $T=64670 2575 0 0 $X=64275 $Y=2235
X65 VDD 21 6 VDD pch_CDNS_764966941092 $T=64670 9755 0 0 $X=64275 $Y=9415
X66 VSS 11 7 VSS nch_CDNS_764966941093 $T=51680 -22660 0 0 $X=51375 $Y=-23000
X67 11 8 9 VSS nch_CDNS_764966941093 $T=51680 -17980 0 0 $X=51375 $Y=-18320
X68 VSS 14 7 VSS nch_CDNS_764966941093 $T=54970 -22660 0 0 $X=54665 $Y=-23000
X69 14 12 8 VSS nch_CDNS_764966941093 $T=54970 -17980 0 0 $X=54665 $Y=-18320
X70 VSS 17 7 VSS nch_CDNS_764966941093 $T=58260 -22660 0 0 $X=57955 $Y=-23000
X71 17 15 12 VSS nch_CDNS_764966941093 $T=58260 -17980 0 0 $X=57955 $Y=-18320
X72 VSS 20 7 VSS nch_CDNS_764966941093 $T=61550 -22660 0 0 $X=61245 $Y=-23000
X73 20 18 15 VSS nch_CDNS_764966941093 $T=61550 -17980 0 0 $X=61245 $Y=-18320
X74 VSS 22 7 VSS nch_CDNS_764966941093 $T=64840 -22660 0 0 $X=64535 $Y=-23000
X75 22 9 18 VSS nch_CDNS_764966941093 $T=64840 -17980 0 0 $X=64535 $Y=-18320
X76 VDD pch_lvt_CDNS_764966941098 $T=77005 -5445 0 0 $X=76610 $Y=-5785
X77 VDD pch_lvt_CDNS_764966941098 $T=77005 1995 0 0 $X=76610 $Y=1655
X78 VDD pch_lvt_CDNS_764966941098 $T=77005 9435 0 0 $X=76610 $Y=9095
X79 VDD pch_lvt_CDNS_764966941098 $T=77005 16875 0 0 $X=76610 $Y=16535
X80 VDD pch_lvt_CDNS_764966941098 $T=82395 -5445 0 0 $X=82000 $Y=-5785
X81 VDD pch_lvt_CDNS_764966941098 $T=82395 16875 0 0 $X=82000 $Y=16535
X82 VDD pch_lvt_CDNS_764966941098 $T=87785 -5445 0 0 $X=87390 $Y=-5785
X83 VDD pch_lvt_CDNS_764966941098 $T=87785 16875 0 0 $X=87390 $Y=16535
X84 VDD pch_lvt_CDNS_764966941098 $T=93175 -5445 0 0 $X=92780 $Y=-5785
X85 VDD pch_lvt_CDNS_764966941098 $T=93175 1995 0 0 $X=92780 $Y=1655
X86 VDD pch_lvt_CDNS_764966941098 $T=93175 9435 0 0 $X=92780 $Y=9095
X87 VDD pch_lvt_CDNS_764966941098 $T=93175 16875 0 0 $X=92780 $Y=16535
X88 VSS nch_lvt_CDNS_764966941099 $T=77020 -34340 0 0 $X=76715 $Y=-34680
X89 VSS nch_lvt_CDNS_764966941099 $T=77020 -27860 0 0 $X=76715 $Y=-28200
X90 VSS nch_lvt_CDNS_764966941099 $T=77020 -21380 0 0 $X=76715 $Y=-21720
X91 VSS nch_lvt_CDNS_764966941099 $T=77020 -14900 0 0 $X=76715 $Y=-15240
X92 VSS nch_lvt_CDNS_764966941099 $T=82410 -34340 0 0 $X=82105 $Y=-34680
X93 VSS nch_lvt_CDNS_764966941099 $T=82410 -14900 0 0 $X=82105 $Y=-15240
X94 VSS nch_lvt_CDNS_764966941099 $T=87800 -34340 0 0 $X=87495 $Y=-34680
X95 VSS nch_lvt_CDNS_764966941099 $T=87800 -14900 0 0 $X=87495 $Y=-15240
X96 VSS nch_lvt_CDNS_764966941099 $T=93190 -34340 0 0 $X=92885 $Y=-34680
X97 VSS nch_lvt_CDNS_764966941099 $T=93190 -27860 0 0 $X=92885 $Y=-28200
X98 VSS nch_lvt_CDNS_764966941099 $T=93190 -21380 0 0 $X=92885 $Y=-21720
X99 VSS nch_lvt_CDNS_764966941099 $T=93190 -14900 0 0 $X=92885 $Y=-15240
X100 VDD 23 9 pch_lvt_CDNS_7649669410913 $T=82395 1995 0 0 $X=82000 $Y=1655
X101 VDD 23 9 pch_lvt_CDNS_7649669410913 $T=82395 9435 0 0 $X=82000 $Y=9095
X102 VDD f_out 23 pch_lvt_CDNS_7649669410913 $T=87785 1995 0 0 $X=87390 $Y=1655
X103 VDD f_out 23 pch_lvt_CDNS_7649669410913 $T=87785 9435 0 0 $X=87390 $Y=9095
X104 VSS 23 9 nch_lvt_CDNS_7649669410910 $T=82410 -27860 0 0 $X=82105 $Y=-28200
X105 VSS 23 9 nch_lvt_CDNS_7649669410910 $T=82410 -21380 0 0 $X=82105 $Y=-21720
X106 VSS f_out 23 nch_lvt_CDNS_7649669410910 $T=87800 -27860 0 0 $X=87495 $Y=-28200
X107 VSS f_out 23 nch_lvt_CDNS_7649669410910 $T=87800 -21380 0 0 $X=87495 $Y=-21720
.ENDS
***************************************
.SUBCKT INVD0BWP7T I VSS VDD ZN
** N=4 EP=4 IP=0 FDC=2
M0 ZN I VSS VSS nch L=6e-08 W=1.5e-07 $X=325 $Y=200 $D=4
M1 ZN I VDD VDD pch L=6e-08 W=1.9e-07 $X=325 $Y=1010 $D=103
.ENDS
***************************************
.SUBCKT ND2D0BWP7T A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=4
M0 6 A2 VSS VSS nch L=6e-08 W=1.5e-07 $X=240 $Y=200 $D=4
M1 ZN A1 6 VSS nch L=6e-08 W=1.5e-07 $X=445 $Y=200 $D=4
M2 ZN A2 VDD VDD pch L=6e-08 W=1.9e-07 $X=240 $Y=1010 $D=103
M3 VDD A1 ZN VDD pch L=6e-08 W=1.9e-07 $X=500 $Y=1010 $D=103
.ENDS
***************************************
.SUBCKT INVD2BWP7T I ZN VDD VSS
** N=4 EP=4 IP=0 FDC=4
M0 ZN I VSS VSS nch L=6e-08 W=3e-07 $X=240 $Y=200 $D=4
M1 VSS I ZN VSS nch L=6e-08 W=3e-07 $X=510 $Y=200 $D=4
M2 ZN I VDD VDD pch L=6e-08 W=3.8e-07 $X=240 $Y=820 $D=103
M3 VDD I ZN VDD pch L=6e-08 W=3.8e-07 $X=510 $Y=820 $D=103
.ENDS
***************************************
.SUBCKT ND3D0BWP7T A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS nch L=6e-08 W=1.5e-07 $X=245 $Y=200 $D=4
M1 8 A2 7 VSS nch L=6e-08 W=1.5e-07 $X=465 $Y=200 $D=4
M2 ZN A1 8 VSS nch L=6e-08 W=1.5e-07 $X=685 $Y=200 $D=4
M3 ZN A3 VDD VDD pch L=6e-08 W=1.9e-07 $X=215 $Y=990 $D=103
M4 VDD A2 ZN VDD pch L=6e-08 W=1.9e-07 $X=475 $Y=990 $D=103
M5 ZN A1 VDD VDD pch L=6e-08 W=1.9e-07 $X=725 $Y=820 $D=103
.ENDS
***************************************
.SUBCKT BUFFD0BWP7T I VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS I 5 VSS nch L=6e-08 W=1.5e-07 $X=225 $Y=200 $D=4
M1 Z 5 VSS VSS nch L=6e-08 W=1.5e-07 $X=505 $Y=200 $D=4
M2 VDD I 5 VDD pch L=6e-08 W=1.9e-07 $X=225 $Y=960 $D=103
M3 Z 5 VDD VDD pch L=6e-08 W=1.9e-07 $X=505 $Y=960 $D=103
.ENDS
***************************************
.SUBCKT PFD BPSK_REG BPSK VDD VSS DN_PFD UP_PFD N_off_PFD P_on_PFD
** N=30 EP=8 IP=98 FDC=84
M0 28 12 VSS VSS nch L=6e-08 W=1.5e-07 $X=6670 $Y=5250 $D=4
M1 29 14 28 VSS nch L=6e-08 W=1.5e-07 $X=6930 $Y=5250 $D=4
M2 30 18 29 VSS nch L=6e-08 W=1.5e-07 $X=7190 $Y=5250 $D=4
M3 13 16 30 VSS nch L=6e-08 W=1.5e-07 $X=7450 $Y=5250 $D=4
M4 13 12 VDD VDD pch L=6e-08 W=1.9e-07 $X=6670 $Y=6060 $D=103
M5 VDD 14 13 VDD pch L=6e-08 W=1.9e-07 $X=6930 $Y=6060 $D=103
M6 13 18 VDD VDD pch L=6e-08 W=1.9e-07 $X=7190 $Y=6060 $D=103
M7 VDD 16 13 VDD pch L=6e-08 W=1.9e-07 $X=7450 $Y=6060 $D=103
X8 BPSK_REG VSS VDD 10 INVD0BWP7T $T=3730 2250 1 0 $X=3495 $Y=615
X9 BPSK VSS VDD 11 INVD0BWP7T $T=3730 7850 0 0 $X=3495 $Y=7745
X10 15 VSS VDD 24 INVD0BWP7T $T=10730 2250 1 0 $X=10495 $Y=615
X11 15 VSS VDD 25 INVD0BWP7T $T=10730 2250 0 0 $X=10495 $Y=2145
X12 19 VSS VDD 26 INVD0BWP7T $T=10730 7850 1 0 $X=10495 $Y=6215
X13 19 VSS VDD 27 INVD0BWP7T $T=10730 7850 0 0 $X=10495 $Y=7745
X14 25 VSS VDD N_off_PFD INVD0BWP7T $T=12130 2250 0 0 $X=11895 $Y=2145
X15 26 VSS VDD P_on_PFD INVD0BWP7T $T=12130 7850 1 0 $X=11895 $Y=6215
X16 15 VSS 10 14 VDD ND2D0BWP7T $T=4930 2250 1 0 $X=4695 $Y=615
X17 14 VSS 17 12 VDD ND2D0BWP7T $T=4930 2250 0 0 $X=4695 $Y=2145
X18 12 VSS 13 17 VDD ND2D0BWP7T $T=4930 5050 1 0 $X=4695 $Y=3415
X19 13 VSS 16 9 VDD ND2D0BWP7T $T=4930 5050 0 0 $X=4695 $Y=4945
X20 9 VSS 18 16 VDD ND2D0BWP7T $T=4930 7850 1 0 $X=4695 $Y=6215
X21 11 VSS 19 18 VDD ND2D0BWP7T $T=4930 7850 0 0 $X=4695 $Y=7745
X22 14 21 VDD VSS INVD2BWP7T $T=6330 2250 1 0 $X=6095 $Y=615
X23 18 20 VDD VSS INVD2BWP7T $T=6330 7850 0 0 $X=6095 $Y=7745
X24 21 23 VDD VSS INVD2BWP7T $T=7730 2250 1 0 $X=7495 $Y=615
X25 20 22 VDD VSS INVD2BWP7T $T=7730 7850 0 0 $X=7495 $Y=7745
X26 23 VSS 12 13 VDD 15 ND3D0BWP7T $T=9130 2250 1 0 $X=8895 $Y=615
X27 13 VSS 16 22 VDD 19 ND3D0BWP7T $T=9130 7850 0 0 $X=8895 $Y=7745
X28 24 VSS VDD DN_PFD BUFFD0BWP7T $T=11930 2250 1 0 $X=11695 $Y=615
X29 27 VSS VDD UP_PFD BUFFD0BWP7T $T=11930 7850 0 0 $X=11695 $Y=7745
.ENDS
***************************************
.SUBCKT pch_lvt_CDNS_7649669410932 1
** N=2 EP=1 IP=0 FDC=1
M0 1 1 1 1 pch_lvt L=1.2e-06 W=3e-07 $X=0 $Y=0 $D=121
.ENDS
***************************************
.SUBCKT ICV_29 1
** N=2 EP=1 IP=4 FDC=2
X0 1 pch_lvt_CDNS_7649669410932 $T=0 0 0 0 $X=-395 $Y=-340
X1 1 pch_lvt_CDNS_7649669410932 $T=0 1160 0 0 $X=-395 $Y=820
.ENDS
***************************************
.SUBCKT ICV_30 1
** N=2 EP=1 IP=4 FDC=4
X0 1 ICV_29 $T=0 0 0 0 $X=-395 $Y=-340
X1 1 ICV_29 $T=0 2320 0 0 $X=-395 $Y=1980
.ENDS
***************************************
.SUBCKT pch_lvt_CDNS_7649669410934 1
** N=2 EP=1 IP=0 FDC=1
M0 1 1 1 1 pch_lvt L=1.2e-06 W=3e-07 $X=0 $Y=0 $D=121
.ENDS
***************************************
.SUBCKT ICV_27 1
** N=2 EP=1 IP=4 FDC=2
X0 1 pch_lvt_CDNS_7649669410934 $T=0 0 0 0 $X=-395 $Y=-340
X1 1 pch_lvt_CDNS_7649669410934 $T=0 1160 0 0 $X=-395 $Y=820
.ENDS
***************************************
.SUBCKT ICV_28 1
** N=2 EP=1 IP=4 FDC=4
X0 1 ICV_27 $T=0 0 0 0 $X=-395 $Y=-340
X1 1 ICV_27 $T=0 2320 0 0 $X=-395 $Y=1980
.ENDS
***************************************
.SUBCKT M1_PO_CDNS_7649669410948
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pch_lvt_CDNS_7649669410929 1 2 3 5
** N=5 EP=4 IP=0 FDC=1
M0 2 3 1 5 pch_lvt L=1.2e-06 W=3e-07 $X=0 $Y=0 $D=121
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 8
** N=8 EP=7 IP=10 FDC=2
X0 1 2 5 8 pch_lvt_CDNS_7649669410929 $T=0 0 0 0 $X=-395 $Y=-340
X1 3 4 6 8 pch_lvt_CDNS_7649669410929 $T=3190 0 1 180 $X=1595 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6 7 9
** N=9 EP=8 IP=16 FDC=4
X0 1 2 4 3 2 6 9 ICV_32 $T=0 0 0 0 $X=-395 $Y=-340
X1 4 5 1 2 7 2 9 ICV_32 $T=0 1160 0 0 $X=-395 $Y=820
.ENDS
***************************************
.SUBCKT ICV_31
** N=3 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT nch_lvt_CDNS_7649669410925 1
** N=1 EP=1 IP=0 FDC=1
M0 1 1 1 1 nch_lvt L=1.2e-06 W=3e-07 $X=0 $Y=0 $D=45
.ENDS
***************************************
.SUBCKT ICV_26 1
** N=1 EP=1 IP=2 FDC=2
X0 1 nch_lvt_CDNS_7649669410925 $T=0 0 0 0 $X=-305 $Y=-340
X1 1 nch_lvt_CDNS_7649669410925 $T=0 1160 0 0 $X=-305 $Y=820
.ENDS
***************************************
.SUBCKT nch_lvt_CDNS_7649669410926 1
** N=1 EP=1 IP=0 FDC=1
M0 1 1 1 1 nch_lvt L=1.2e-06 W=1.2e-06 $X=0 $Y=0 $D=45
.ENDS
***************************************
.SUBCKT pch_lvt_CDNS_7649669410931 1
** N=2 EP=1 IP=0 FDC=1
M0 1 1 1 1 pch_lvt L=1.2e-06 W=1.2e-06 $X=0 $Y=0 $D=121
.ENDS
***************************************
.SUBCKT nch_lvt_CDNS_7649669410928 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch_lvt L=1.2e-06 W=3e-07 $X=0 $Y=0 $D=45
.ENDS
***************************************
.SUBCKT nch_lvt_CDNS_7649669410927 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nch_lvt L=1.2e-06 W=1.2e-06 $X=0 $Y=0 $D=45
.ENDS
***************************************
.SUBCKT pch_lvt_CDNS_7649669410930 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch_lvt L=1.2e-06 W=1.2e-06 $X=0 $Y=0 $D=121
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410935 1
** N=1 EP=1 IP=0 FDC=1
M0 1 1 1 1 nch L=3e-07 W=3e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_24 1
** N=1 EP=1 IP=2 FDC=2
X0 1 nch_CDNS_7649669410935 $T=0 0 0 0 $X=-305 $Y=-340
X1 1 nch_CDNS_7649669410935 $T=1025 0 0 0 $X=720 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_25 1
** N=1 EP=1 IP=2 FDC=4
X0 1 ICV_24 $T=0 0 0 0 $X=-305 $Y=-340
X1 1 ICV_24 $T=2050 0 0 0 $X=1745 $Y=-340
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410923 1
** N=1 EP=1 IP=0 FDC=1
M0 1 1 1 1 nch L=6e-08 W=1.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT pch_CDNS_7649669410924 1
** N=2 EP=1 IP=0 FDC=1
M0 1 1 1 1 pch L=6e-08 W=2.4e-07 $X=0 $Y=0 $D=103
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410916 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=3e-07 W=3e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3
** N=3 EP=3 IP=6 FDC=2
X0 1 2 3 nch_CDNS_7649669410916 $T=0 0 0 0 $X=-305 $Y=-340
X1 1 2 3 nch_CDNS_7649669410916 $T=1025 0 0 0 $X=720 $Y=-340
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410920 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nch L=6e-08 W=1.2e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT pch_CDNS_7649669410921 1 2 3 5
** N=5 EP=4 IP=0 FDC=1
M0 2 3 1 5 pch L=6e-08 W=2.4e-07 $X=0 $Y=0 $D=103
.ENDS
***************************************
.SUBCKT nch_CDNS_7649669410917 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nch L=3e-07 W=3e-07 $X=0 $Y=0 $D=4
.ENDS
***************************************
.SUBCKT pch_CDNS_7649669410922 1
** N=2 EP=1 IP=0 FDC=1
M0 1 1 1 1 pch L=3e-07 W=6e-07 $X=0 $Y=0 $D=103
.ENDS
***************************************
.SUBCKT ICV_21 1
** N=2 EP=1 IP=4 FDC=2
X0 1 pch_CDNS_7649669410922 $T=0 0 0 0 $X=-395 $Y=-340
X1 1 pch_CDNS_7649669410922 $T=1090 0 0 0 $X=695 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_20 1
** N=2 EP=1 IP=4 FDC=2
X0 1 pch_CDNS_7649669410922 $T=0 0 0 0 $X=-395 $Y=-340
X1 1 pch_CDNS_7649669410922 $T=0 1460 0 0 $X=-395 $Y=1120
.ENDS
***************************************
.SUBCKT pch_CDNS_7649669410919 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pch L=3e-07 W=6e-07 $X=0 $Y=0 $D=103
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3
** N=4 EP=3 IP=8 FDC=2
X0 1 2 3 pch_CDNS_7649669410919 $T=0 0 0 0 $X=-395 $Y=-340
X1 1 2 3 pch_CDNS_7649669410919 $T=1090 0 0 0 $X=695 $Y=-340
.ENDS
***************************************
.SUBCKT Charge_pump VDD GND CP_out CR_1uA_CP_OP CR_1uA_CP N_off_CP P_on_CP UP_CP DN_CP
** N=19 EP=9 IP=601 FDC=278
M0 19 19 VDD VDD pch L=3e-07 W=6e-07 $X=97090 $Y=51660 $D=103
X1 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=61650 $Y=29900 $D=325
X2 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=61650 $Y=41300 $D=325
X3 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=61650 $Y=52700 $D=325
X4 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=69850 $Y=29900 $D=325
X5 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=69850 $Y=41300 $D=325
X6 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=69850 $Y=52700 $D=325
X7 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=78050 $Y=29900 $D=325
X8 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=78050 $Y=41300 $D=325
X9 13 14 mimcap_sin lt=4e-06 wt=4e-06 mimflag=3 $X=78050 $Y=52700 $D=325
X10 VDD pch_lvt_CDNS_7649669410932 $T=65160 13480 0 0 $X=64765 $Y=13140
X11 VDD pch_lvt_CDNS_7649669410932 $T=65160 23920 0 0 $X=64765 $Y=23580
X12 VDD pch_lvt_CDNS_7649669410932 $T=67150 13480 0 0 $X=66755 $Y=13140
X13 VDD pch_lvt_CDNS_7649669410932 $T=67150 23920 0 0 $X=66755 $Y=23580
X14 VDD ICV_29 $T=63170 22760 0 0 $X=62775 $Y=22420
X15 VDD ICV_29 $T=69140 22760 0 0 $X=68745 $Y=22420
X16 VDD ICV_30 $T=63170 13480 0 0 $X=62775 $Y=13140
X17 VDD ICV_30 $T=63170 18120 0 0 $X=62775 $Y=17780
X18 VDD ICV_30 $T=69140 13480 0 0 $X=68745 $Y=13140
X19 VDD ICV_30 $T=69140 18120 0 0 $X=68745 $Y=17780
X20 VDD pch_lvt_CDNS_7649669410934 $T=63170 39340 0 0 $X=62775 $Y=39000
X21 VDD pch_lvt_CDNS_7649669410934 $T=65160 27740 0 0 $X=64765 $Y=27400
X22 VDD pch_lvt_CDNS_7649669410934 $T=65160 39340 0 0 $X=64765 $Y=39000
X23 VDD pch_lvt_CDNS_7649669410934 $T=67150 27740 0 0 $X=66755 $Y=27400
X24 VDD pch_lvt_CDNS_7649669410934 $T=67150 39340 0 0 $X=66755 $Y=39000
X25 VDD pch_lvt_CDNS_7649669410934 $T=69140 39340 0 0 $X=68745 $Y=39000
X26 VDD ICV_27 $T=63170 37020 0 0 $X=62775 $Y=36680
X27 VDD ICV_27 $T=69140 37020 0 0 $X=68745 $Y=36680
X28 VDD ICV_28 $T=63170 27740 0 0 $X=62775 $Y=27400
X29 VDD ICV_28 $T=63170 32380 0 0 $X=62775 $Y=32040
X30 VDD ICV_28 $T=69140 27740 0 0 $X=68745 $Y=27400
X31 VDD ICV_28 $T=69140 32380 0 0 $X=68745 $Y=32040
X96 VDD 10 VDD 14 10 11 VDD ICV_32 $T=65160 38180 0 0 $X=64765 $Y=37840
X97 10 12 13 11 13 12 12 VDD ICV_33 $T=65160 14640 0 0 $X=64765 $Y=14300
X98 10 12 13 11 13 12 12 VDD ICV_33 $T=65160 16960 0 0 $X=64765 $Y=16620
X99 10 12 13 11 13 12 12 VDD ICV_33 $T=65160 19280 0 0 $X=64765 $Y=18940
X100 10 12 13 11 13 12 12 VDD ICV_33 $T=65160 21600 0 0 $X=64765 $Y=21260
X101 VDD 10 10 VDD 14 10 11 VDD ICV_33 $T=65160 28900 0 0 $X=64765 $Y=28560
X102 VDD 10 14 VDD 14 11 11 VDD ICV_33 $T=65160 31220 0 0 $X=64765 $Y=30880
X103 VDD 10 14 VDD 14 11 11 VDD ICV_33 $T=65160 33540 0 0 $X=64765 $Y=33200
X104 VDD 10 14 VDD 14 11 11 VDD ICV_33 $T=65160 35860 0 0 $X=64765 $Y=35520
X118 GND nch_lvt_CDNS_7649669410925 $T=75790 13310 0 0 $X=75485 $Y=12970
X119 GND nch_lvt_CDNS_7649669410925 $T=75790 19110 0 0 $X=75485 $Y=18770
X120 GND nch_lvt_CDNS_7649669410925 $T=77780 13310 0 0 $X=77475 $Y=12970
X121 GND nch_lvt_CDNS_7649669410925 $T=77780 19110 0 0 $X=77475 $Y=18770
X122 GND ICV_26 $T=73800 13310 0 0 $X=73495 $Y=12970
X123 GND ICV_26 $T=73800 15630 0 0 $X=73495 $Y=15290
X124 GND ICV_26 $T=73800 17950 0 0 $X=73495 $Y=17610
X125 GND ICV_26 $T=79770 13310 0 0 $X=79465 $Y=12970
X126 GND ICV_26 $T=79770 15630 0 0 $X=79465 $Y=15290
X127 GND ICV_26 $T=79770 17950 0 0 $X=79465 $Y=17610
X128 GND nch_lvt_CDNS_7649669410926 $T=73800 22590 0 0 $X=73495 $Y=22250
X129 GND nch_lvt_CDNS_7649669410926 $T=73800 24650 0 0 $X=73495 $Y=24310
X130 GND nch_lvt_CDNS_7649669410926 $T=73800 26710 0 0 $X=73495 $Y=26370
X131 GND nch_lvt_CDNS_7649669410926 $T=73800 28770 0 0 $X=73495 $Y=28430
X132 GND nch_lvt_CDNS_7649669410926 $T=75790 22590 0 0 $X=75485 $Y=22250
X133 GND nch_lvt_CDNS_7649669410926 $T=75790 28770 0 0 $X=75485 $Y=28430
X134 GND nch_lvt_CDNS_7649669410926 $T=77780 22590 0 0 $X=77475 $Y=22250
X135 GND nch_lvt_CDNS_7649669410926 $T=77780 28770 0 0 $X=77475 $Y=28430
X136 GND nch_lvt_CDNS_7649669410926 $T=79770 22590 0 0 $X=79465 $Y=22250
X137 GND nch_lvt_CDNS_7649669410926 $T=79770 24650 0 0 $X=79465 $Y=24310
X138 GND nch_lvt_CDNS_7649669410926 $T=79770 26710 0 0 $X=79465 $Y=26370
X139 GND nch_lvt_CDNS_7649669410926 $T=79770 28770 0 0 $X=79465 $Y=28430
X140 VDD pch_lvt_CDNS_7649669410931 $T=73970 33320 0 0 $X=73575 $Y=32980
X141 VDD pch_lvt_CDNS_7649669410931 $T=73970 35380 0 0 $X=73575 $Y=35040
X142 VDD pch_lvt_CDNS_7649669410931 $T=73970 37440 0 0 $X=73575 $Y=37100
X143 VDD pch_lvt_CDNS_7649669410931 $T=73970 39500 0 0 $X=73575 $Y=39160
X144 VDD pch_lvt_CDNS_7649669410931 $T=75960 33320 0 0 $X=75565 $Y=32980
X145 VDD pch_lvt_CDNS_7649669410931 $T=75960 39500 0 0 $X=75565 $Y=39160
X146 VDD pch_lvt_CDNS_7649669410931 $T=77950 33320 0 0 $X=77555 $Y=32980
X147 VDD pch_lvt_CDNS_7649669410931 $T=77950 39500 0 0 $X=77555 $Y=39160
X148 VDD pch_lvt_CDNS_7649669410931 $T=79940 33320 0 0 $X=79545 $Y=32980
X149 VDD pch_lvt_CDNS_7649669410931 $T=79940 35380 0 0 $X=79545 $Y=35040
X150 VDD pch_lvt_CDNS_7649669410931 $T=79940 37440 0 0 $X=79545 $Y=37100
X151 VDD pch_lvt_CDNS_7649669410931 $T=79940 39500 0 0 $X=79545 $Y=39160
X152 GND CR_1uA_CP_OP CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=75790 14470 0 0 $X=75485 $Y=14130
X153 GND 14 CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=75790 15630 0 0 $X=75485 $Y=15290
X154 GND 12 CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=75790 16790 0 0 $X=75485 $Y=16450
X155 GND 15 CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=75790 17950 0 0 $X=75485 $Y=17610
X156 GND 15 CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=78980 14470 1 180 $X=77475 $Y=14130
X157 GND 12 CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=78980 15630 1 180 $X=77475 $Y=15290
X158 GND 14 CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=78980 16790 1 180 $X=77475 $Y=16450
X159 GND CR_1uA_CP_OP CR_1uA_CP_OP nch_lvt_CDNS_7649669410928 $T=78980 17950 1 180 $X=77475 $Y=17610
X160 15 11 CP_out GND nch_lvt_CDNS_7649669410927 $T=75790 24650 0 0 $X=75485 $Y=24310
X161 15 16 14 GND nch_lvt_CDNS_7649669410927 $T=75790 26710 0 0 $X=75485 $Y=26370
X162 15 16 14 GND nch_lvt_CDNS_7649669410927 $T=78980 24650 1 180 $X=77475 $Y=24310
X163 15 11 CP_out GND nch_lvt_CDNS_7649669410927 $T=78980 26710 1 180 $X=77475 $Y=26370
X164 VDD 11 16 pch_lvt_CDNS_7649669410930 $T=75960 35380 0 0 $X=75565 $Y=35040
X165 VDD 16 16 pch_lvt_CDNS_7649669410930 $T=75960 37440 0 0 $X=75565 $Y=37100
X166 VDD 16 16 pch_lvt_CDNS_7649669410930 $T=79150 35380 1 180 $X=77555 $Y=35040
X167 VDD 11 16 pch_lvt_CDNS_7649669410930 $T=79150 37440 1 180 $X=77555 $Y=37100
X168 GND nch_CDNS_7649669410935 $T=87130 39850 0 0 $X=86825 $Y=39510
X169 GND nch_CDNS_7649669410935 $T=87130 41010 0 0 $X=86825 $Y=40670
X170 GND nch_CDNS_7649669410935 $T=99430 38690 0 0 $X=99125 $Y=38350
X171 GND nch_CDNS_7649669410935 $T=99430 39850 0 0 $X=99125 $Y=39510
X172 GND nch_CDNS_7649669410935 $T=99430 41010 0 0 $X=99125 $Y=40670
X173 GND nch_CDNS_7649669410935 $T=99430 42170 0 0 $X=99125 $Y=41830
X174 GND ICV_25 $T=87130 38690 0 0 $X=86825 $Y=38350
X175 GND ICV_25 $T=87130 42170 0 0 $X=86825 $Y=41830
X176 GND ICV_25 $T=91230 38690 0 0 $X=90925 $Y=38350
X177 GND ICV_25 $T=91230 42170 0 0 $X=90925 $Y=41830
X178 GND ICV_25 $T=95330 38690 0 0 $X=95025 $Y=38350
X179 GND ICV_25 $T=95330 42170 0 0 $X=95025 $Y=41830
X180 GND nch_CDNS_7649669410923 $T=87640 45660 0 0 $X=87260 $Y=45320
X181 GND nch_CDNS_7649669410923 $T=87640 46640 0 0 $X=87260 $Y=46300
X182 GND nch_CDNS_7649669410923 $T=87640 47620 0 0 $X=87260 $Y=47280
X183 GND nch_CDNS_7649669410923 $T=87640 48600 0 0 $X=87260 $Y=48260
X184 GND nch_CDNS_7649669410923 $T=88640 45660 0 0 $X=88260 $Y=45320
X185 GND nch_CDNS_7649669410923 $T=88640 48600 0 0 $X=88260 $Y=48260
X186 GND nch_CDNS_7649669410923 $T=89640 45660 0 0 $X=89260 $Y=45320
X187 GND nch_CDNS_7649669410923 $T=89640 48600 0 0 $X=89260 $Y=48260
X188 GND nch_CDNS_7649669410923 $T=90640 45660 0 0 $X=90260 $Y=45320
X189 GND nch_CDNS_7649669410923 $T=90640 46640 0 0 $X=90260 $Y=46300
X190 GND nch_CDNS_7649669410923 $T=90640 47620 0 0 $X=90260 $Y=47280
X191 GND nch_CDNS_7649669410923 $T=90640 48600 0 0 $X=90260 $Y=48260
X192 VDD pch_CDNS_7649669410924 $T=87865 54060 0 0 $X=87470 $Y=53720
X193 VDD pch_CDNS_7649669410924 $T=87865 55160 0 0 $X=87470 $Y=54820
X194 VDD pch_CDNS_7649669410924 $T=87865 56260 0 0 $X=87470 $Y=55920
X195 VDD pch_CDNS_7649669410924 $T=87865 57360 0 0 $X=87470 $Y=57020
X196 VDD pch_CDNS_7649669410924 $T=88715 54060 0 0 $X=88320 $Y=53720
X197 VDD pch_CDNS_7649669410924 $T=88715 57360 0 0 $X=88320 $Y=57020
X198 VDD pch_CDNS_7649669410924 $T=89565 54060 0 0 $X=89170 $Y=53720
X199 VDD pch_CDNS_7649669410924 $T=89565 57360 0 0 $X=89170 $Y=57020
X200 VDD pch_CDNS_7649669410924 $T=90415 54060 0 0 $X=90020 $Y=53720
X201 VDD pch_CDNS_7649669410924 $T=90415 55160 0 0 $X=90020 $Y=54820
X202 VDD pch_CDNS_7649669410924 $T=90415 56260 0 0 $X=90020 $Y=55920
X203 VDD pch_CDNS_7649669410924 $T=90415 57360 0 0 $X=90020 $Y=57020
X204 GND 17 CR_1uA_CP nch_CDNS_7649669410916 $T=92255 39850 0 0 $X=91950 $Y=39510
X205 GND 17 CR_1uA_CP nch_CDNS_7649669410916 $T=92255 41010 0 0 $X=91950 $Y=40670
X206 GND 17 CR_1uA_CP nch_CDNS_7649669410916 $T=98405 39850 0 0 $X=98100 $Y=39510
X207 GND 17 CR_1uA_CP nch_CDNS_7649669410916 $T=98405 41010 0 0 $X=98100 $Y=40670
X208 GND 17 CR_1uA_CP ICV_22 $T=88155 39850 0 0 $X=87850 $Y=39510
X209 GND 17 CR_1uA_CP ICV_22 $T=88155 41010 0 0 $X=87850 $Y=40670
X210 GND 17 CR_1uA_CP ICV_22 $T=90205 39850 0 0 $X=89900 $Y=39510
X211 GND 17 CR_1uA_CP ICV_22 $T=90205 41010 0 0 $X=89900 $Y=40670
X212 GND 17 CR_1uA_CP ICV_22 $T=94305 39850 0 0 $X=94000 $Y=39510
X213 GND 17 CR_1uA_CP ICV_22 $T=94305 41010 0 0 $X=94000 $Y=40670
X214 GND 17 CR_1uA_CP ICV_22 $T=96355 39850 0 0 $X=96050 $Y=39510
X215 GND 17 CR_1uA_CP ICV_22 $T=96355 41010 0 0 $X=96050 $Y=40670
X216 17 14 N_off_CP GND nch_CDNS_7649669410920 $T=88640 46640 0 0 $X=88260 $Y=46300
X217 17 CP_out DN_CP GND nch_CDNS_7649669410920 $T=88640 47620 0 0 $X=88260 $Y=47280
X218 17 CP_out DN_CP GND nch_CDNS_7649669410920 $T=89700 46640 1 180 $X=89260 $Y=46300
X219 17 14 N_off_CP GND nch_CDNS_7649669410920 $T=89700 47620 1 180 $X=89260 $Y=47280
X220 18 CP_out P_on_CP VDD pch_CDNS_7649669410921 $T=88715 55160 0 0 $X=88320 $Y=54820
X221 18 14 UP_CP VDD pch_CDNS_7649669410921 $T=88715 56260 0 0 $X=88320 $Y=55920
X222 18 14 UP_CP VDD pch_CDNS_7649669410921 $T=89625 55160 1 180 $X=89170 $Y=54820
X223 18 CP_out P_on_CP VDD pch_CDNS_7649669410921 $T=89625 56260 1 180 $X=89170 $Y=55920
X224 GND CR_1uA_CP CR_1uA_CP nch_CDNS_7649669410917 $T=93280 39850 0 0 $X=92975 $Y=39510
X225 GND 19 CR_1uA_CP nch_CDNS_7649669410917 $T=93280 41010 0 0 $X=92975 $Y=40670
X226 VDD pch_CDNS_7649669410922 $T=94910 56040 0 0 $X=94515 $Y=55700
X227 VDD pch_CDNS_7649669410922 $T=99270 57500 0 0 $X=98875 $Y=57160
X228 VDD ICV_21 $T=94910 45820 0 0 $X=94515 $Y=45480
X229 VDD ICV_21 $T=94910 57500 0 0 $X=94515 $Y=57160
X230 VDD ICV_21 $T=97090 45820 0 0 $X=96695 $Y=45480
X231 VDD ICV_21 $T=97090 57500 0 0 $X=96695 $Y=57160
X232 VDD ICV_20 $T=94910 47280 0 0 $X=94515 $Y=46940
X233 VDD ICV_20 $T=94910 50200 0 0 $X=94515 $Y=49860
X234 VDD ICV_20 $T=94910 53120 0 0 $X=94515 $Y=52780
X235 VDD ICV_20 $T=99270 45820 0 0 $X=98875 $Y=45480
X236 VDD ICV_20 $T=99270 48740 0 0 $X=98875 $Y=48400
X237 VDD ICV_20 $T=99270 51660 0 0 $X=98875 $Y=51320
X238 VDD ICV_20 $T=99270 54580 0 0 $X=98875 $Y=54240
X239 VDD 18 19 pch_CDNS_7649669410919 $T=96000 51660 0 0 $X=95605 $Y=51320
X240 VDD 18 19 pch_CDNS_7649669410919 $T=98180 47280 0 0 $X=97785 $Y=46940
X241 VDD 18 19 pch_CDNS_7649669410919 $T=98180 48740 0 0 $X=97785 $Y=48400
X242 VDD 18 19 pch_CDNS_7649669410919 $T=98180 50200 0 0 $X=97785 $Y=49860
X243 VDD 18 19 pch_CDNS_7649669410919 $T=98180 51660 0 0 $X=97785 $Y=51320
X244 VDD 18 19 pch_CDNS_7649669410919 $T=98180 53120 0 0 $X=97785 $Y=52780
X245 VDD 18 19 pch_CDNS_7649669410919 $T=98180 54580 0 0 $X=97785 $Y=54240
X246 VDD 18 19 pch_CDNS_7649669410919 $T=98180 56040 0 0 $X=97785 $Y=55700
X247 VDD 18 19 ICV_23 $T=96000 47280 0 0 $X=95605 $Y=46940
X248 VDD 18 19 ICV_23 $T=96000 48740 0 0 $X=95605 $Y=48400
X249 VDD 18 19 ICV_23 $T=96000 50200 0 0 $X=95605 $Y=49860
X250 VDD 18 19 ICV_23 $T=96000 53120 0 0 $X=95605 $Y=52780
X251 VDD 18 19 ICV_23 $T=96000 54580 0 0 $X=95605 $Y=54240
X252 VDD 18 19 ICV_23 $T=96000 56040 0 0 $X=95605 $Y=55700
.ENDS
***************************************
.SUBCKT PLL_25M_400M VDD VSS CP_20u_Bias CP_OP_1u_bias f_out input_clk div_sel[0] div_sel[1] div_sel[2] div_sel[3] reset DVDD
** N=19 EP=12 IP=40 FDC=3139
X0 1 3 rppolywo l=1.2e-05 w=2e-06 $X=228675 $Y=-276815 $D=486
X1 1 VSS mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=29905 $Y=-331650 $D=325
X2 1 VSS mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=88265 $Y=-391250 $D=325
X3 1 VSS mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=88265 $Y=-331650 $D=325
X4 1 VSS mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=146625 $Y=-391250 $D=325
X5 1 VSS mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=146625 $Y=-331650 $D=325
X6 1 VSS mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=204985 $Y=-391250 $D=325
X7 1 VSS mimcap_sin lt=5e-05 wt=5e-05 mimflag=3 $X=204985 $Y=-331650 $D=325
X8 VSS 1 mimcap_CDNS_764966941090 $T=29905 -391250 0 0 $X=19505 $Y=-403650
X9 VSS 1 mimcap_CDNS_764966941090 $T=29905 -272050 0 0 $X=19505 $Y=-284450
X10 VSS 1 mimcap_CDNS_764966941090 $T=88265 -272050 0 0 $X=77865 $Y=-284450
X11 VSS 1 mimcap_CDNS_764966941090 $T=263345 -391250 0 0 $X=252945 $Y=-403650
X12 VSS 3 mimcap_CDNS_764966941090 $T=263345 -331650 0 0 $X=252945 $Y=-344050
X13 DVDD VSS 8 f_out reset div_sel[1] div_sel[2] div_sel[3] div_sel[0] clk_div $T=193665 -279650 0 90 $X=151765 $Y=-277150
X14 3 VDD VSS f_out Ring_VCO $T=297490 -234645 1 180 $X=200050 $Y=-270625
X15 8 input_clk VDD VSS 12 11 13 10 PFD $T=253740 -221225 0 0 $X=256135 $Y=-221110
X16 VDD VSS 3 CP_20u_Bias CP_OP_1u_bias 13 10 11 12 Charge_pump $T=374995 -278750 1 180 $X=274210 $Y=-266430
.ENDS
***************************************
